// ============================================================================
// Project:   SPHINCSLET
// Description:   Keccak Round Module
//
//
// This code is almost a straight translation of the VHDL high-speed module
// provided from http://keccak.noekeon.org/.
//
// The MIT License (MIT)
//
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
// ============================================================================


module keccak_round 
#(
    parameter N = 64
)
(
    input   [1599:0]        Round_in,
    input   [N-1:0]         Round_constant_signal,
    output  [1599:0]        Round_out
    );


wire [N-1:0] theta_in [4:0][4:0];
wire [N-1:0] theta_out[4:0][4:0];
wire [N-1:0] pi_in    [4:0][4:0];
wire [N-1:0] pi_out   [4:0][4:0];
wire [N-1:0] rho_in   [4:0][4:0];
wire [N-1:0] rho_out  [4:0][4:0];
wire [N-1:0] chi_in   [4:0][4:0];
wire [N-1:0] chi_out  [4:0][4:0];
wire [N-1:0] iota_in  [4:0][4:0];
wire [N-1:0] iota_out [4:0][4:0];


// k_plane sum_sheet;

wire [N-1:0] sum_sheet[4:0];

wire [N-1:0] round_in_map [4:0][4:0];
wire [N-1:0] round_out_map[4:0][4:0];


genvar i,j,k;
generate        
    for(i=0; i<5; i=i+1) begin
        for (j=0; j<5; j=j+1) begin
            for (k=0; k<64; k=k+1) begin
                assign round_in_map[i][j][k] = Round_in[64*(24-(5*i+j))+k];
            end
        end
    end
endgenerate

// Function: k_state to bit array
generate
    for(i=0; i<5; i=i+1) begin
        for (j=0; j<5; j=j+1) begin
            for (k=0; k<64; k=k+1) begin
                assign Round_out[64*(24-(5*i+j))+k] = round_out_map[i][j][k];
            end
        end
    end
endgenerate


// Connections

// Order is theta, pi, rho, chi, iota
genvar i_i, j_j;
generate
    for (i_i = 0; i_i < 5; i_i = i_i + 1) begin
        for (j_j = 0; j_j < 5; j_j = j_j + 1) begin
            assign  theta_in[i_i][j_j]          = round_in_map[i_i][j_j];
            assign  pi_in[i_i][j_j]             = rho_out[i_i][j_j];
            assign  rho_in[i_i][j_j]            = theta_out[i_i][j_j];
            assign  chi_in[i_i][j_j]            = pi_out[i_i][j_j];
            assign  iota_in[i_i][j_j]           = chi_out[i_i][j_j];
            assign  round_out_map[i_i][j_j]     = iota_out[i_i][j_j];
        end
    end
endgenerate




// Chi
genvar y, x, z;
generate
    for (y = 0; y <= 4; y = y + 1) begin
        for (x = 0; x <= 2; x = x + 1) begin
            for (z = 0; z <= N-1; z = z + 1) begin
                assign chi_out[y][x][z] = chi_in[y][x][z] ^ (~(chi_in[y][x+1][z]) & chi_in[y][x+2][z]);
            end
        end
    end
endgenerate


genvar yy, ii;
generate
    for (yy = 0; yy <= 4; yy = yy + 1) begin
        for (ii = 0; ii <= N-1; ii = ii + 1) begin
            assign chi_out[yy][3][ii] = chi_in[yy][3][ii] ^ (~(chi_in[yy][4][ii]) & chi_in[yy][0][ii]);
        end
    end
endgenerate


genvar yyy, iii;
generate
   for (yyy = 0; yyy <= 4; yyy = yyy+ 1) begin 
       for (iii = 0; iii <= N-1; iii = iii + 1) begin 
           assign chi_out[yyy][4][iii] = chi_in[yyy][4][iii] ^ (~(chi_in[yyy][0][iii]) & chi_in[yyy][1][iii]);
       end
   end
endgenerate



genvar xx, jj;
generate
    for (xx = 0; xx <= 4; xx = xx + 1) begin 
        for (jj = 0; jj <= N-1; jj = jj + 1) begin 
            assign sum_sheet[xx][jj] = theta_in[0][xx][jj] ^ theta_in[1][xx][jj] ^ theta_in[2][xx][jj] ^ theta_in[3][xx][jj] ^ theta_in[4][xx][jj];
        end
    end
endgenerate


genvar m,n,o;
generate
    for(m = 0; m <= 4; m = m + 1) begin 
        for(n = 1; n <= 3; n = n + 1) begin
            assign theta_out[m][n][0] = theta_in[m][n][0] ^ sum_sheet[n-1][0] ^ sum_sheet[n+1][N-1];

            for(o = 1; o <= N-1; o = o + 1) begin 
                assign theta_out[m][n][o] = theta_in[m][n][o] ^ sum_sheet[n-1][o] ^ sum_sheet[n+1][o-1];
            end
        end
    end
endgenerate



genvar mm, oo;
generate
    for(mm = 0; mm <= 4; mm = mm + 1) begin
        assign theta_out[mm][0][0] = theta_in[mm][0][0] ^ sum_sheet[4][0] ^ sum_sheet[1][N-1];

        for(oo = 1; oo <= N-1; oo = oo + 1) begin 
            assign theta_out[mm][0][oo] = theta_in[mm][0][oo] ^ sum_sheet[4][oo] ^ sum_sheet[1][oo-1];
        end
    end
endgenerate


genvar p, q;
generate
    for(p = 0; p <= 4; p = p + 1) begin 
        assign theta_out[p][4][0] = theta_in[p][4][0] ^ sum_sheet[3][0] ^ sum_sheet[0][N-1];

        for(q = 1; q <= N-1; q = q + 1) begin 
            assign theta_out[p][4][q] = theta_in[p][4][q] ^ sum_sheet[3][q] ^ sum_sheet[0][q-1];
        end
    end
endgenerate


genvar pp,qq,rr;
generate
    for (pp = 0; pp <= 4; pp = pp + 1) begin
        for (qq = 0; qq <= 4; qq = qq + 1) begin
            for (rr = 0; rr <= N-1; rr = rr + 1) begin
                assign pi_out[(2*qq+3*pp) % 5][0*qq+1*pp][rr] = pi_in[pp][qq][rr];
            end
        end
    end
endgenerate



genvar f, g, h;
generate
    for (f = 1; f <= 4; f = f + 1) begin 
        for (g = 0; g <= 4; g = g + 1) begin
            for (h = 0; h <= N-1; h = h + 1) begin
                assign iota_out[f][g][h] = iota_in[f][g][h];
            end
        end
    end
endgenerate


genvar ff, gg;
generate
    for (ff = 1; ff <= 4; ff = ff + 1) begin 
        for (gg = 0; gg <= N-1; gg = gg + 1) begin 
            assign iota_out[0][ff][gg] = iota_in[0][ff][gg];
        end
    end
endgenerate


assign rho_out[0][0][ 0 ] = rho_in[0][0][ 0 ];
assign rho_out[0][1][ 0 ] = rho_in[0][1][ 63 ];
assign rho_out[0][2][ 0 ] = rho_in[0][2][ 2 ];
assign rho_out[0][3][ 0 ] = rho_in[0][3][ 36 ];
assign rho_out[0][4][ 0 ] = rho_in[0][4][ 37 ];
assign rho_out[1][0][ 0 ] = rho_in[1][0][ 28 ];
assign rho_out[1][1][ 0 ] = rho_in[1][1][ 20 ];
assign rho_out[1][2][ 0 ] = rho_in[1][2][ 58 ];
assign rho_out[1][3][ 0 ] = rho_in[1][3][ 9 ];
assign rho_out[1][4][ 0 ] = rho_in[1][4][ 44 ];
assign rho_out[2][0][ 0 ] = rho_in[2][0][ 61 ];
assign rho_out[2][1][ 0 ] = rho_in[2][1][ 54 ];
assign rho_out[2][2][ 0 ] = rho_in[2][2][ 21 ];
assign rho_out[2][3][ 0 ] = rho_in[2][3][ 39 ];
assign rho_out[2][4][ 0 ] = rho_in[2][4][ 25 ];
assign rho_out[3][0][ 0 ] = rho_in[3][0][ 23 ];
assign rho_out[3][1][ 0 ] = rho_in[3][1][ 19 ];
assign rho_out[3][2][ 0 ] = rho_in[3][2][ 49 ];
assign rho_out[3][3][ 0 ] = rho_in[3][3][ 43 ];
assign rho_out[3][4][ 0 ] = rho_in[3][4][ 56 ];
assign rho_out[4][0][ 0 ] = rho_in[4][0][ 46 ];
assign rho_out[4][1][ 0 ] = rho_in[4][1][ 62 ];
assign rho_out[4][2][ 0 ] = rho_in[4][2][ 3 ];
assign rho_out[4][3][ 0 ] = rho_in[4][3][ 8 ];
assign rho_out[4][4][ 0 ] = rho_in[4][4][ 50 ];
assign rho_out[0][0][ 1 ] = rho_in[0][0][ 1 ];
assign rho_out[0][1][ 1 ] = rho_in[0][1][ 0 ];
assign rho_out[0][2][ 1 ] = rho_in[0][2][ 3 ];
assign rho_out[0][3][ 1 ] = rho_in[0][3][ 37 ];
assign rho_out[0][4][ 1 ] = rho_in[0][4][ 38 ];
assign rho_out[1][0][ 1 ] = rho_in[1][0][ 29 ];
assign rho_out[1][1][ 1 ] = rho_in[1][1][ 21 ];
assign rho_out[1][2][ 1 ] = rho_in[1][2][ 59 ];
assign rho_out[1][3][ 1 ] = rho_in[1][3][ 10 ];
assign rho_out[1][4][ 1 ] = rho_in[1][4][ 45 ];
assign rho_out[2][0][ 1 ] = rho_in[2][0][ 62 ];
assign rho_out[2][1][ 1 ] = rho_in[2][1][ 55 ];
assign rho_out[2][2][ 1 ] = rho_in[2][2][ 22 ];
assign rho_out[2][3][ 1 ] = rho_in[2][3][ 40 ];
assign rho_out[2][4][ 1 ] = rho_in[2][4][ 26 ];
assign rho_out[3][0][ 1 ] = rho_in[3][0][ 24 ];
assign rho_out[3][1][ 1 ] = rho_in[3][1][ 20 ];
assign rho_out[3][2][ 1 ] = rho_in[3][2][ 50 ];
assign rho_out[3][3][ 1 ] = rho_in[3][3][ 44 ];
assign rho_out[3][4][ 1 ] = rho_in[3][4][ 57 ];
assign rho_out[4][0][ 1 ] = rho_in[4][0][ 47 ];
assign rho_out[4][1][ 1 ] = rho_in[4][1][ 63 ];
assign rho_out[4][2][ 1 ] = rho_in[4][2][ 4 ];
assign rho_out[4][3][ 1 ] = rho_in[4][3][ 9 ];
assign rho_out[4][4][ 1 ] = rho_in[4][4][ 51 ];
assign rho_out[0][0][ 2 ] = rho_in[0][0][ 2 ];
assign rho_out[0][1][ 2 ] = rho_in[0][1][ 1 ];
assign rho_out[0][2][ 2 ] = rho_in[0][2][ 4 ];
assign rho_out[0][3][ 2 ] = rho_in[0][3][ 38 ];
assign rho_out[0][4][ 2 ] = rho_in[0][4][ 39 ];
assign rho_out[1][0][ 2 ] = rho_in[1][0][ 30 ];
assign rho_out[1][1][ 2 ] = rho_in[1][1][ 22 ];
assign rho_out[1][2][ 2 ] = rho_in[1][2][ 60 ];
assign rho_out[1][3][ 2 ] = rho_in[1][3][ 11 ];
assign rho_out[1][4][ 2 ] = rho_in[1][4][ 46 ];
assign rho_out[2][0][ 2 ] = rho_in[2][0][ 63 ];
assign rho_out[2][1][ 2 ] = rho_in[2][1][ 56 ];
assign rho_out[2][2][ 2 ] = rho_in[2][2][ 23 ];
assign rho_out[2][3][ 2 ] = rho_in[2][3][ 41 ];
assign rho_out[2][4][ 2 ] = rho_in[2][4][ 27 ];
assign rho_out[3][0][ 2 ] = rho_in[3][0][ 25 ];
assign rho_out[3][1][ 2 ] = rho_in[3][1][ 21 ];
assign rho_out[3][2][ 2 ] = rho_in[3][2][ 51 ];
assign rho_out[3][3][ 2 ] = rho_in[3][3][ 45 ];
assign rho_out[3][4][ 2 ] = rho_in[3][4][ 58 ];
assign rho_out[4][0][ 2 ] = rho_in[4][0][ 48 ];
assign rho_out[4][1][ 2 ] = rho_in[4][1][ 0 ];
assign rho_out[4][2][ 2 ] = rho_in[4][2][ 5 ];
assign rho_out[4][3][ 2 ] = rho_in[4][3][ 10 ];
assign rho_out[4][4][ 2 ] = rho_in[4][4][ 52 ];
assign rho_out[0][0][ 3 ] = rho_in[0][0][ 3 ];
assign rho_out[0][1][ 3 ] = rho_in[0][1][ 2 ];
assign rho_out[0][2][ 3 ] = rho_in[0][2][ 5 ];
assign rho_out[0][3][ 3 ] = rho_in[0][3][ 39 ];
assign rho_out[0][4][ 3 ] = rho_in[0][4][ 40 ];
assign rho_out[1][0][ 3 ] = rho_in[1][0][ 31 ];
assign rho_out[1][1][ 3 ] = rho_in[1][1][ 23 ];
assign rho_out[1][2][ 3 ] = rho_in[1][2][ 61 ];
assign rho_out[1][3][ 3 ] = rho_in[1][3][ 12 ];
assign rho_out[1][4][ 3 ] = rho_in[1][4][ 47 ];
assign rho_out[2][0][ 3 ] = rho_in[2][0][ 0 ];
assign rho_out[2][1][ 3 ] = rho_in[2][1][ 57 ];
assign rho_out[2][2][ 3 ] = rho_in[2][2][ 24 ];
assign rho_out[2][3][ 3 ] = rho_in[2][3][ 42 ];
assign rho_out[2][4][ 3 ] = rho_in[2][4][ 28 ];
assign rho_out[3][0][ 3 ] = rho_in[3][0][ 26 ];
assign rho_out[3][1][ 3 ] = rho_in[3][1][ 22 ];
assign rho_out[3][2][ 3 ] = rho_in[3][2][ 52 ];
assign rho_out[3][3][ 3 ] = rho_in[3][3][ 46 ];
assign rho_out[3][4][ 3 ] = rho_in[3][4][ 59 ];
assign rho_out[4][0][ 3 ] = rho_in[4][0][ 49 ];
assign rho_out[4][1][ 3 ] = rho_in[4][1][ 1 ];
assign rho_out[4][2][ 3 ] = rho_in[4][2][ 6 ];
assign rho_out[4][3][ 3 ] = rho_in[4][3][ 11 ];
assign rho_out[4][4][ 3 ] = rho_in[4][4][ 53 ];
assign rho_out[0][0][ 4 ] = rho_in[0][0][ 4 ];
assign rho_out[0][1][ 4 ] = rho_in[0][1][ 3 ];
assign rho_out[0][2][ 4 ] = rho_in[0][2][ 6 ];
assign rho_out[0][3][ 4 ] = rho_in[0][3][ 40 ];
assign rho_out[0][4][ 4 ] = rho_in[0][4][ 41 ];
assign rho_out[1][0][ 4 ] = rho_in[1][0][ 32 ];
assign rho_out[1][1][ 4 ] = rho_in[1][1][ 24 ];
assign rho_out[1][2][ 4 ] = rho_in[1][2][ 62 ];
assign rho_out[1][3][ 4 ] = rho_in[1][3][ 13 ];
assign rho_out[1][4][ 4 ] = rho_in[1][4][ 48 ];
assign rho_out[2][0][ 4 ] = rho_in[2][0][ 1 ];
assign rho_out[2][1][ 4 ] = rho_in[2][1][ 58 ];
assign rho_out[2][2][ 4 ] = rho_in[2][2][ 25 ];
assign rho_out[2][3][ 4 ] = rho_in[2][3][ 43 ];
assign rho_out[2][4][ 4 ] = rho_in[2][4][ 29 ];
assign rho_out[3][0][ 4 ] = rho_in[3][0][ 27 ];
assign rho_out[3][1][ 4 ] = rho_in[3][1][ 23 ];
assign rho_out[3][2][ 4 ] = rho_in[3][2][ 53 ];
assign rho_out[3][3][ 4 ] = rho_in[3][3][ 47 ];
assign rho_out[3][4][ 4 ] = rho_in[3][4][ 60 ];
assign rho_out[4][0][ 4 ] = rho_in[4][0][ 50 ];
assign rho_out[4][1][ 4 ] = rho_in[4][1][ 2 ];
assign rho_out[4][2][ 4 ] = rho_in[4][2][ 7 ];
assign rho_out[4][3][ 4 ] = rho_in[4][3][ 12 ];
assign rho_out[4][4][ 4 ] = rho_in[4][4][ 54 ];
assign rho_out[0][0][ 5 ] = rho_in[0][0][ 5 ];
assign rho_out[0][1][ 5 ] = rho_in[0][1][ 4 ];
assign rho_out[0][2][ 5 ] = rho_in[0][2][ 7 ];
assign rho_out[0][3][ 5 ] = rho_in[0][3][ 41 ];
assign rho_out[0][4][ 5 ] = rho_in[0][4][ 42 ];
assign rho_out[1][0][ 5 ] = rho_in[1][0][ 33 ];
assign rho_out[1][1][ 5 ] = rho_in[1][1][ 25 ];
assign rho_out[1][2][ 5 ] = rho_in[1][2][ 63 ];
assign rho_out[1][3][ 5 ] = rho_in[1][3][ 14 ];
assign rho_out[1][4][ 5 ] = rho_in[1][4][ 49 ];
assign rho_out[2][0][ 5 ] = rho_in[2][0][ 2 ];
assign rho_out[2][1][ 5 ] = rho_in[2][1][ 59 ];
assign rho_out[2][2][ 5 ] = rho_in[2][2][ 26 ];
assign rho_out[2][3][ 5 ] = rho_in[2][3][ 44 ];
assign rho_out[2][4][ 5 ] = rho_in[2][4][ 30 ];
assign rho_out[3][0][ 5 ] = rho_in[3][0][ 28 ];
assign rho_out[3][1][ 5 ] = rho_in[3][1][ 24 ];
assign rho_out[3][2][ 5 ] = rho_in[3][2][ 54 ];
assign rho_out[3][3][ 5 ] = rho_in[3][3][ 48 ];
assign rho_out[3][4][ 5 ] = rho_in[3][4][ 61 ];
assign rho_out[4][0][ 5 ] = rho_in[4][0][ 51 ];
assign rho_out[4][1][ 5 ] = rho_in[4][1][ 3 ];
assign rho_out[4][2][ 5 ] = rho_in[4][2][ 8 ];
assign rho_out[4][3][ 5 ] = rho_in[4][3][ 13 ];
assign rho_out[4][4][ 5 ] = rho_in[4][4][ 55 ];
assign rho_out[0][0][ 6 ] = rho_in[0][0][ 6 ];
assign rho_out[0][1][ 6 ] = rho_in[0][1][ 5 ];
assign rho_out[0][2][ 6 ] = rho_in[0][2][ 8 ];
assign rho_out[0][3][ 6 ] = rho_in[0][3][ 42 ];
assign rho_out[0][4][ 6 ] = rho_in[0][4][ 43 ];
assign rho_out[1][0][ 6 ] = rho_in[1][0][ 34 ];
assign rho_out[1][1][ 6 ] = rho_in[1][1][ 26 ];
assign rho_out[1][2][ 6 ] = rho_in[1][2][ 0 ];
assign rho_out[1][3][ 6 ] = rho_in[1][3][ 15 ];
assign rho_out[1][4][ 6 ] = rho_in[1][4][ 50 ];
assign rho_out[2][0][ 6 ] = rho_in[2][0][ 3 ];
assign rho_out[2][1][ 6 ] = rho_in[2][1][ 60 ];
assign rho_out[2][2][ 6 ] = rho_in[2][2][ 27 ];
assign rho_out[2][3][ 6 ] = rho_in[2][3][ 45 ];
assign rho_out[2][4][ 6 ] = rho_in[2][4][ 31 ];
assign rho_out[3][0][ 6 ] = rho_in[3][0][ 29 ];
assign rho_out[3][1][ 6 ] = rho_in[3][1][ 25 ];
assign rho_out[3][2][ 6 ] = rho_in[3][2][ 55 ];
assign rho_out[3][3][ 6 ] = rho_in[3][3][ 49 ];
assign rho_out[3][4][ 6 ] = rho_in[3][4][ 62 ];
assign rho_out[4][0][ 6 ] = rho_in[4][0][ 52 ];
assign rho_out[4][1][ 6 ] = rho_in[4][1][ 4 ];
assign rho_out[4][2][ 6 ] = rho_in[4][2][ 9 ];
assign rho_out[4][3][ 6 ] = rho_in[4][3][ 14 ];
assign rho_out[4][4][ 6 ] = rho_in[4][4][ 56 ];
assign rho_out[0][0][ 7 ] = rho_in[0][0][ 7 ];
assign rho_out[0][1][ 7 ] = rho_in[0][1][ 6 ];
assign rho_out[0][2][ 7 ] = rho_in[0][2][ 9 ];
assign rho_out[0][3][ 7 ] = rho_in[0][3][ 43 ];
assign rho_out[0][4][ 7 ] = rho_in[0][4][ 44 ];
assign rho_out[1][0][ 7 ] = rho_in[1][0][ 35 ];
assign rho_out[1][1][ 7 ] = rho_in[1][1][ 27 ];
assign rho_out[1][2][ 7 ] = rho_in[1][2][ 1 ];
assign rho_out[1][3][ 7 ] = rho_in[1][3][ 16 ];
assign rho_out[1][4][ 7 ] = rho_in[1][4][ 51 ];
assign rho_out[2][0][ 7 ] = rho_in[2][0][ 4 ];
assign rho_out[2][1][ 7 ] = rho_in[2][1][ 61 ];
assign rho_out[2][2][ 7 ] = rho_in[2][2][ 28 ];
assign rho_out[2][3][ 7 ] = rho_in[2][3][ 46 ];
assign rho_out[2][4][ 7 ] = rho_in[2][4][ 32 ];
assign rho_out[3][0][ 7 ] = rho_in[3][0][ 30 ];
assign rho_out[3][1][ 7 ] = rho_in[3][1][ 26 ];
assign rho_out[3][2][ 7 ] = rho_in[3][2][ 56 ];
assign rho_out[3][3][ 7 ] = rho_in[3][3][ 50 ];
assign rho_out[3][4][ 7 ] = rho_in[3][4][ 63 ];
assign rho_out[4][0][ 7 ] = rho_in[4][0][ 53 ];
assign rho_out[4][1][ 7 ] = rho_in[4][1][ 5 ];
assign rho_out[4][2][ 7 ] = rho_in[4][2][ 10 ];
assign rho_out[4][3][ 7 ] = rho_in[4][3][ 15 ];
assign rho_out[4][4][ 7 ] = rho_in[4][4][ 57 ];
assign rho_out[0][0][ 8 ] = rho_in[0][0][ 8 ];
assign rho_out[0][1][ 8 ] = rho_in[0][1][ 7 ];
assign rho_out[0][2][ 8 ] = rho_in[0][2][ 10 ];
assign rho_out[0][3][ 8 ] = rho_in[0][3][ 44 ];
assign rho_out[0][4][ 8 ] = rho_in[0][4][ 45 ];
assign rho_out[1][0][ 8 ] = rho_in[1][0][ 36 ];
assign rho_out[1][1][ 8 ] = rho_in[1][1][ 28 ];
assign rho_out[1][2][ 8 ] = rho_in[1][2][ 2 ];
assign rho_out[1][3][ 8 ] = rho_in[1][3][ 17 ];
assign rho_out[1][4][ 8 ] = rho_in[1][4][ 52 ];
assign rho_out[2][0][ 8 ] = rho_in[2][0][ 5 ];
assign rho_out[2][1][ 8 ] = rho_in[2][1][ 62 ];
assign rho_out[2][2][ 8 ] = rho_in[2][2][ 29 ];
assign rho_out[2][3][ 8 ] = rho_in[2][3][ 47 ];
assign rho_out[2][4][ 8 ] = rho_in[2][4][ 33 ];
assign rho_out[3][0][ 8 ] = rho_in[3][0][ 31 ];
assign rho_out[3][1][ 8 ] = rho_in[3][1][ 27 ];
assign rho_out[3][2][ 8 ] = rho_in[3][2][ 57 ];
assign rho_out[3][3][ 8 ] = rho_in[3][3][ 51 ];
assign rho_out[3][4][ 8 ] = rho_in[3][4][ 0 ];
assign rho_out[4][0][ 8 ] = rho_in[4][0][ 54 ];
assign rho_out[4][1][ 8 ] = rho_in[4][1][ 6 ];
assign rho_out[4][2][ 8 ] = rho_in[4][2][ 11 ];
assign rho_out[4][3][ 8 ] = rho_in[4][3][ 16 ];
assign rho_out[4][4][ 8 ] = rho_in[4][4][ 58 ];
assign rho_out[0][0][ 9 ] = rho_in[0][0][ 9 ];
assign rho_out[0][1][ 9 ] = rho_in[0][1][ 8 ];
assign rho_out[0][2][ 9 ] = rho_in[0][2][ 11 ];
assign rho_out[0][3][ 9 ] = rho_in[0][3][ 45 ];
assign rho_out[0][4][ 9 ] = rho_in[0][4][ 46 ];
assign rho_out[1][0][ 9 ] = rho_in[1][0][ 37 ];
assign rho_out[1][1][ 9 ] = rho_in[1][1][ 29 ];
assign rho_out[1][2][ 9 ] = rho_in[1][2][ 3 ];
assign rho_out[1][3][ 9 ] = rho_in[1][3][ 18 ];
assign rho_out[1][4][ 9 ] = rho_in[1][4][ 53 ];
assign rho_out[2][0][ 9 ] = rho_in[2][0][ 6 ];
assign rho_out[2][1][ 9 ] = rho_in[2][1][ 63 ];
assign rho_out[2][2][ 9 ] = rho_in[2][2][ 30 ];
assign rho_out[2][3][ 9 ] = rho_in[2][3][ 48 ];
assign rho_out[2][4][ 9 ] = rho_in[2][4][ 34 ];
assign rho_out[3][0][ 9 ] = rho_in[3][0][ 32 ];
assign rho_out[3][1][ 9 ] = rho_in[3][1][ 28 ];
assign rho_out[3][2][ 9 ] = rho_in[3][2][ 58 ];
assign rho_out[3][3][ 9 ] = rho_in[3][3][ 52 ];
assign rho_out[3][4][ 9 ] = rho_in[3][4][ 1 ];
assign rho_out[4][0][ 9 ] = rho_in[4][0][ 55 ];
assign rho_out[4][1][ 9 ] = rho_in[4][1][ 7 ];
assign rho_out[4][2][ 9 ] = rho_in[4][2][ 12 ];
assign rho_out[4][3][ 9 ] = rho_in[4][3][ 17 ];
assign rho_out[4][4][ 9 ] = rho_in[4][4][ 59 ];
assign rho_out[0][0][ 10 ] = rho_in[0][0][ 10 ];
assign rho_out[0][1][ 10 ] = rho_in[0][1][ 9 ];
assign rho_out[0][2][ 10 ] = rho_in[0][2][ 12 ];
assign rho_out[0][3][ 10 ] = rho_in[0][3][ 46 ];
assign rho_out[0][4][ 10 ] = rho_in[0][4][ 47 ];
assign rho_out[1][0][ 10 ] = rho_in[1][0][ 38 ];
assign rho_out[1][1][ 10 ] = rho_in[1][1][ 30 ];
assign rho_out[1][2][ 10 ] = rho_in[1][2][ 4 ];
assign rho_out[1][3][ 10 ] = rho_in[1][3][ 19 ];
assign rho_out[1][4][ 10 ] = rho_in[1][4][ 54 ];
assign rho_out[2][0][ 10 ] = rho_in[2][0][ 7 ];
assign rho_out[2][1][ 10 ] = rho_in[2][1][ 0 ];
assign rho_out[2][2][ 10 ] = rho_in[2][2][ 31 ];
assign rho_out[2][3][ 10 ] = rho_in[2][3][ 49 ];
assign rho_out[2][4][ 10 ] = rho_in[2][4][ 35 ];
assign rho_out[3][0][ 10 ] = rho_in[3][0][ 33 ];
assign rho_out[3][1][ 10 ] = rho_in[3][1][ 29 ];
assign rho_out[3][2][ 10 ] = rho_in[3][2][ 59 ];
assign rho_out[3][3][ 10 ] = rho_in[3][3][ 53 ];
assign rho_out[3][4][ 10 ] = rho_in[3][4][ 2 ];
assign rho_out[4][0][ 10 ] = rho_in[4][0][ 56 ];
assign rho_out[4][1][ 10 ] = rho_in[4][1][ 8 ];
assign rho_out[4][2][ 10 ] = rho_in[4][2][ 13 ];
assign rho_out[4][3][ 10 ] = rho_in[4][3][ 18 ];
assign rho_out[4][4][ 10 ] = rho_in[4][4][ 60 ];
assign rho_out[0][0][ 11 ] = rho_in[0][0][ 11 ];
assign rho_out[0][1][ 11 ] = rho_in[0][1][ 10 ];
assign rho_out[0][2][ 11 ] = rho_in[0][2][ 13 ];
assign rho_out[0][3][ 11 ] = rho_in[0][3][ 47 ];
assign rho_out[0][4][ 11 ] = rho_in[0][4][ 48 ];
assign rho_out[1][0][ 11 ] = rho_in[1][0][ 39 ];
assign rho_out[1][1][ 11 ] = rho_in[1][1][ 31 ];
assign rho_out[1][2][ 11 ] = rho_in[1][2][ 5 ];
assign rho_out[1][3][ 11 ] = rho_in[1][3][ 20 ];
assign rho_out[1][4][ 11 ] = rho_in[1][4][ 55 ];
assign rho_out[2][0][ 11 ] = rho_in[2][0][ 8 ];
assign rho_out[2][1][ 11 ] = rho_in[2][1][ 1 ];
assign rho_out[2][2][ 11 ] = rho_in[2][2][ 32 ];
assign rho_out[2][3][ 11 ] = rho_in[2][3][ 50 ];
assign rho_out[2][4][ 11 ] = rho_in[2][4][ 36 ];
assign rho_out[3][0][ 11 ] = rho_in[3][0][ 34 ];
assign rho_out[3][1][ 11 ] = rho_in[3][1][ 30 ];
assign rho_out[3][2][ 11 ] = rho_in[3][2][ 60 ];
assign rho_out[3][3][ 11 ] = rho_in[3][3][ 54 ];
assign rho_out[3][4][ 11 ] = rho_in[3][4][ 3 ];
assign rho_out[4][0][ 11 ] = rho_in[4][0][ 57 ];
assign rho_out[4][1][ 11 ] = rho_in[4][1][ 9 ];
assign rho_out[4][2][ 11 ] = rho_in[4][2][ 14 ];
assign rho_out[4][3][ 11 ] = rho_in[4][3][ 19 ];
assign rho_out[4][4][ 11 ] = rho_in[4][4][ 61 ];
assign rho_out[0][0][ 12 ] = rho_in[0][0][ 12 ];
assign rho_out[0][1][ 12 ] = rho_in[0][1][ 11 ];
assign rho_out[0][2][ 12 ] = rho_in[0][2][ 14 ];
assign rho_out[0][3][ 12 ] = rho_in[0][3][ 48 ];
assign rho_out[0][4][ 12 ] = rho_in[0][4][ 49 ];
assign rho_out[1][0][ 12 ] = rho_in[1][0][ 40 ];
assign rho_out[1][1][ 12 ] = rho_in[1][1][ 32 ];
assign rho_out[1][2][ 12 ] = rho_in[1][2][ 6 ];
assign rho_out[1][3][ 12 ] = rho_in[1][3][ 21 ];
assign rho_out[1][4][ 12 ] = rho_in[1][4][ 56 ];
assign rho_out[2][0][ 12 ] = rho_in[2][0][ 9 ];
assign rho_out[2][1][ 12 ] = rho_in[2][1][ 2 ];
assign rho_out[2][2][ 12 ] = rho_in[2][2][ 33 ];
assign rho_out[2][3][ 12 ] = rho_in[2][3][ 51 ];
assign rho_out[2][4][ 12 ] = rho_in[2][4][ 37 ];
assign rho_out[3][0][ 12 ] = rho_in[3][0][ 35 ];
assign rho_out[3][1][ 12 ] = rho_in[3][1][ 31 ];
assign rho_out[3][2][ 12 ] = rho_in[3][2][ 61 ];
assign rho_out[3][3][ 12 ] = rho_in[3][3][ 55 ];
assign rho_out[3][4][ 12 ] = rho_in[3][4][ 4 ];
assign rho_out[4][0][ 12 ] = rho_in[4][0][ 58 ];
assign rho_out[4][1][ 12 ] = rho_in[4][1][ 10 ];
assign rho_out[4][2][ 12 ] = rho_in[4][2][ 15 ];
assign rho_out[4][3][ 12 ] = rho_in[4][3][ 20 ];
assign rho_out[4][4][ 12 ] = rho_in[4][4][ 62 ];
assign rho_out[0][0][ 13 ] = rho_in[0][0][ 13 ];
assign rho_out[0][1][ 13 ] = rho_in[0][1][ 12 ];
assign rho_out[0][2][ 13 ] = rho_in[0][2][ 15 ];
assign rho_out[0][3][ 13 ] = rho_in[0][3][ 49 ];
assign rho_out[0][4][ 13 ] = rho_in[0][4][ 50 ];
assign rho_out[1][0][ 13 ] = rho_in[1][0][ 41 ];
assign rho_out[1][1][ 13 ] = rho_in[1][1][ 33 ];
assign rho_out[1][2][ 13 ] = rho_in[1][2][ 7 ];
assign rho_out[1][3][ 13 ] = rho_in[1][3][ 22 ];
assign rho_out[1][4][ 13 ] = rho_in[1][4][ 57 ];
assign rho_out[2][0][ 13 ] = rho_in[2][0][ 10 ];
assign rho_out[2][1][ 13 ] = rho_in[2][1][ 3 ];
assign rho_out[2][2][ 13 ] = rho_in[2][2][ 34 ];
assign rho_out[2][3][ 13 ] = rho_in[2][3][ 52 ];
assign rho_out[2][4][ 13 ] = rho_in[2][4][ 38 ];
assign rho_out[3][0][ 13 ] = rho_in[3][0][ 36 ];
assign rho_out[3][1][ 13 ] = rho_in[3][1][ 32 ];
assign rho_out[3][2][ 13 ] = rho_in[3][2][ 62 ];
assign rho_out[3][3][ 13 ] = rho_in[3][3][ 56 ];
assign rho_out[3][4][ 13 ] = rho_in[3][4][ 5 ];
assign rho_out[4][0][ 13 ] = rho_in[4][0][ 59 ];
assign rho_out[4][1][ 13 ] = rho_in[4][1][ 11 ];
assign rho_out[4][2][ 13 ] = rho_in[4][2][ 16 ];
assign rho_out[4][3][ 13 ] = rho_in[4][3][ 21 ];
assign rho_out[4][4][ 13 ] = rho_in[4][4][ 63 ];
assign rho_out[0][0][ 14 ] = rho_in[0][0][ 14 ];
assign rho_out[0][1][ 14 ] = rho_in[0][1][ 13 ];
assign rho_out[0][2][ 14 ] = rho_in[0][2][ 16 ];
assign rho_out[0][3][ 14 ] = rho_in[0][3][ 50 ];
assign rho_out[0][4][ 14 ] = rho_in[0][4][ 51 ];
assign rho_out[1][0][ 14 ] = rho_in[1][0][ 42 ];
assign rho_out[1][1][ 14 ] = rho_in[1][1][ 34 ];
assign rho_out[1][2][ 14 ] = rho_in[1][2][ 8 ];
assign rho_out[1][3][ 14 ] = rho_in[1][3][ 23 ];
assign rho_out[1][4][ 14 ] = rho_in[1][4][ 58 ];
assign rho_out[2][0][ 14 ] = rho_in[2][0][ 11 ];
assign rho_out[2][1][ 14 ] = rho_in[2][1][ 4 ];
assign rho_out[2][2][ 14 ] = rho_in[2][2][ 35 ];
assign rho_out[2][3][ 14 ] = rho_in[2][3][ 53 ];
assign rho_out[2][4][ 14 ] = rho_in[2][4][ 39 ];
assign rho_out[3][0][ 14 ] = rho_in[3][0][ 37 ];
assign rho_out[3][1][ 14 ] = rho_in[3][1][ 33 ];
assign rho_out[3][2][ 14 ] = rho_in[3][2][ 63 ];
assign rho_out[3][3][ 14 ] = rho_in[3][3][ 57 ];
assign rho_out[3][4][ 14 ] = rho_in[3][4][ 6 ];
assign rho_out[4][0][ 14 ] = rho_in[4][0][ 60 ];
assign rho_out[4][1][ 14 ] = rho_in[4][1][ 12 ];
assign rho_out[4][2][ 14 ] = rho_in[4][2][ 17 ];
assign rho_out[4][3][ 14 ] = rho_in[4][3][ 22 ];
assign rho_out[4][4][ 14 ] = rho_in[4][4][ 0 ];
assign rho_out[0][0][ 15 ] = rho_in[0][0][ 15 ];
assign rho_out[0][1][ 15 ] = rho_in[0][1][ 14 ];
assign rho_out[0][2][ 15 ] = rho_in[0][2][ 17 ];
assign rho_out[0][3][ 15 ] = rho_in[0][3][ 51 ];
assign rho_out[0][4][ 15 ] = rho_in[0][4][ 52 ];
assign rho_out[1][0][ 15 ] = rho_in[1][0][ 43 ];
assign rho_out[1][1][ 15 ] = rho_in[1][1][ 35 ];
assign rho_out[1][2][ 15 ] = rho_in[1][2][ 9 ];
assign rho_out[1][3][ 15 ] = rho_in[1][3][ 24 ];
assign rho_out[1][4][ 15 ] = rho_in[1][4][ 59 ];
assign rho_out[2][0][ 15 ] = rho_in[2][0][ 12 ];
assign rho_out[2][1][ 15 ] = rho_in[2][1][ 5 ];
assign rho_out[2][2][ 15 ] = rho_in[2][2][ 36 ];
assign rho_out[2][3][ 15 ] = rho_in[2][3][ 54 ];
assign rho_out[2][4][ 15 ] = rho_in[2][4][ 40 ];
assign rho_out[3][0][ 15 ] = rho_in[3][0][ 38 ];
assign rho_out[3][1][ 15 ] = rho_in[3][1][ 34 ];
assign rho_out[3][2][ 15 ] = rho_in[3][2][ 0 ];
assign rho_out[3][3][ 15 ] = rho_in[3][3][ 58 ];
assign rho_out[3][4][ 15 ] = rho_in[3][4][ 7 ];
assign rho_out[4][0][ 15 ] = rho_in[4][0][ 61 ];
assign rho_out[4][1][ 15 ] = rho_in[4][1][ 13 ];
assign rho_out[4][2][ 15 ] = rho_in[4][2][ 18 ];
assign rho_out[4][3][ 15 ] = rho_in[4][3][ 23 ];
assign rho_out[4][4][ 15 ] = rho_in[4][4][ 1 ];
assign rho_out[0][0][ 16 ] = rho_in[0][0][ 16 ];
assign rho_out[0][1][ 16 ] = rho_in[0][1][ 15 ];
assign rho_out[0][2][ 16 ] = rho_in[0][2][ 18 ];
assign rho_out[0][3][ 16 ] = rho_in[0][3][ 52 ];
assign rho_out[0][4][ 16 ] = rho_in[0][4][ 53 ];
assign rho_out[1][0][ 16 ] = rho_in[1][0][ 44 ];
assign rho_out[1][1][ 16 ] = rho_in[1][1][ 36 ];
assign rho_out[1][2][ 16 ] = rho_in[1][2][ 10 ];
assign rho_out[1][3][ 16 ] = rho_in[1][3][ 25 ];
assign rho_out[1][4][ 16 ] = rho_in[1][4][ 60 ];
assign rho_out[2][0][ 16 ] = rho_in[2][0][ 13 ];
assign rho_out[2][1][ 16 ] = rho_in[2][1][ 6 ];
assign rho_out[2][2][ 16 ] = rho_in[2][2][ 37 ];
assign rho_out[2][3][ 16 ] = rho_in[2][3][ 55 ];
assign rho_out[2][4][ 16 ] = rho_in[2][4][ 41 ];
assign rho_out[3][0][ 16 ] = rho_in[3][0][ 39 ];
assign rho_out[3][1][ 16 ] = rho_in[3][1][ 35 ];
assign rho_out[3][2][ 16 ] = rho_in[3][2][ 1 ];
assign rho_out[3][3][ 16 ] = rho_in[3][3][ 59 ];
assign rho_out[3][4][ 16 ] = rho_in[3][4][ 8 ];
assign rho_out[4][0][ 16 ] = rho_in[4][0][ 62 ];
assign rho_out[4][1][ 16 ] = rho_in[4][1][ 14 ];
assign rho_out[4][2][ 16 ] = rho_in[4][2][ 19 ];
assign rho_out[4][3][ 16 ] = rho_in[4][3][ 24 ];
assign rho_out[4][4][ 16 ] = rho_in[4][4][ 2 ];
assign rho_out[0][0][ 17 ] = rho_in[0][0][ 17 ];
assign rho_out[0][1][ 17 ] = rho_in[0][1][ 16 ];
assign rho_out[0][2][ 17 ] = rho_in[0][2][ 19 ];
assign rho_out[0][3][ 17 ] = rho_in[0][3][ 53 ];
assign rho_out[0][4][ 17 ] = rho_in[0][4][ 54 ];
assign rho_out[1][0][ 17 ] = rho_in[1][0][ 45 ];
assign rho_out[1][1][ 17 ] = rho_in[1][1][ 37 ];
assign rho_out[1][2][ 17 ] = rho_in[1][2][ 11 ];
assign rho_out[1][3][ 17 ] = rho_in[1][3][ 26 ];
assign rho_out[1][4][ 17 ] = rho_in[1][4][ 61 ];
assign rho_out[2][0][ 17 ] = rho_in[2][0][ 14 ];
assign rho_out[2][1][ 17 ] = rho_in[2][1][ 7 ];
assign rho_out[2][2][ 17 ] = rho_in[2][2][ 38 ];
assign rho_out[2][3][ 17 ] = rho_in[2][3][ 56 ];
assign rho_out[2][4][ 17 ] = rho_in[2][4][ 42 ];
assign rho_out[3][0][ 17 ] = rho_in[3][0][ 40 ];
assign rho_out[3][1][ 17 ] = rho_in[3][1][ 36 ];
assign rho_out[3][2][ 17 ] = rho_in[3][2][ 2 ];
assign rho_out[3][3][ 17 ] = rho_in[3][3][ 60 ];
assign rho_out[3][4][ 17 ] = rho_in[3][4][ 9 ];
assign rho_out[4][0][ 17 ] = rho_in[4][0][ 63 ];
assign rho_out[4][1][ 17 ] = rho_in[4][1][ 15 ];
assign rho_out[4][2][ 17 ] = rho_in[4][2][ 20 ];
assign rho_out[4][3][ 17 ] = rho_in[4][3][ 25 ];
assign rho_out[4][4][ 17 ] = rho_in[4][4][ 3 ];
assign rho_out[0][0][ 18 ] = rho_in[0][0][ 18 ];
assign rho_out[0][1][ 18 ] = rho_in[0][1][ 17 ];
assign rho_out[0][2][ 18 ] = rho_in[0][2][ 20 ];
assign rho_out[0][3][ 18 ] = rho_in[0][3][ 54 ];
assign rho_out[0][4][ 18 ] = rho_in[0][4][ 55 ];
assign rho_out[1][0][ 18 ] = rho_in[1][0][ 46 ];
assign rho_out[1][1][ 18 ] = rho_in[1][1][ 38 ];
assign rho_out[1][2][ 18 ] = rho_in[1][2][ 12 ];
assign rho_out[1][3][ 18 ] = rho_in[1][3][ 27 ];
assign rho_out[1][4][ 18 ] = rho_in[1][4][ 62 ];
assign rho_out[2][0][ 18 ] = rho_in[2][0][ 15 ];
assign rho_out[2][1][ 18 ] = rho_in[2][1][ 8 ];
assign rho_out[2][2][ 18 ] = rho_in[2][2][ 39 ];
assign rho_out[2][3][ 18 ] = rho_in[2][3][ 57 ];
assign rho_out[2][4][ 18 ] = rho_in[2][4][ 43 ];
assign rho_out[3][0][ 18 ] = rho_in[3][0][ 41 ];
assign rho_out[3][1][ 18 ] = rho_in[3][1][ 37 ];
assign rho_out[3][2][ 18 ] = rho_in[3][2][ 3 ];
assign rho_out[3][3][ 18 ] = rho_in[3][3][ 61 ];
assign rho_out[3][4][ 18 ] = rho_in[3][4][ 10 ];
assign rho_out[4][0][ 18 ] = rho_in[4][0][ 0 ];
assign rho_out[4][1][ 18 ] = rho_in[4][1][ 16 ];
assign rho_out[4][2][ 18 ] = rho_in[4][2][ 21 ];
assign rho_out[4][3][ 18 ] = rho_in[4][3][ 26 ];
assign rho_out[4][4][ 18 ] = rho_in[4][4][ 4 ];
assign rho_out[0][0][ 19 ] = rho_in[0][0][ 19 ];
assign rho_out[0][1][ 19 ] = rho_in[0][1][ 18 ];
assign rho_out[0][2][ 19 ] = rho_in[0][2][ 21 ];
assign rho_out[0][3][ 19 ] = rho_in[0][3][ 55 ];
assign rho_out[0][4][ 19 ] = rho_in[0][4][ 56 ];
assign rho_out[1][0][ 19 ] = rho_in[1][0][ 47 ];
assign rho_out[1][1][ 19 ] = rho_in[1][1][ 39 ];
assign rho_out[1][2][ 19 ] = rho_in[1][2][ 13 ];
assign rho_out[1][3][ 19 ] = rho_in[1][3][ 28 ];
assign rho_out[1][4][ 19 ] = rho_in[1][4][ 63 ];
assign rho_out[2][0][ 19 ] = rho_in[2][0][ 16 ];
assign rho_out[2][1][ 19 ] = rho_in[2][1][ 9 ];
assign rho_out[2][2][ 19 ] = rho_in[2][2][ 40 ];
assign rho_out[2][3][ 19 ] = rho_in[2][3][ 58 ];
assign rho_out[2][4][ 19 ] = rho_in[2][4][ 44 ];
assign rho_out[3][0][ 19 ] = rho_in[3][0][ 42 ];
assign rho_out[3][1][ 19 ] = rho_in[3][1][ 38 ];
assign rho_out[3][2][ 19 ] = rho_in[3][2][ 4 ];
assign rho_out[3][3][ 19 ] = rho_in[3][3][ 62 ];
assign rho_out[3][4][ 19 ] = rho_in[3][4][ 11 ];
assign rho_out[4][0][ 19 ] = rho_in[4][0][ 1 ];
assign rho_out[4][1][ 19 ] = rho_in[4][1][ 17 ];
assign rho_out[4][2][ 19 ] = rho_in[4][2][ 22 ];
assign rho_out[4][3][ 19 ] = rho_in[4][3][ 27 ];
assign rho_out[4][4][ 19 ] = rho_in[4][4][ 5 ];
assign rho_out[0][0][ 20 ] = rho_in[0][0][ 20 ];
assign rho_out[0][1][ 20 ] = rho_in[0][1][ 19 ];
assign rho_out[0][2][ 20 ] = rho_in[0][2][ 22 ];
assign rho_out[0][3][ 20 ] = rho_in[0][3][ 56 ];
assign rho_out[0][4][ 20 ] = rho_in[0][4][ 57 ];
assign rho_out[1][0][ 20 ] = rho_in[1][0][ 48 ];
assign rho_out[1][1][ 20 ] = rho_in[1][1][ 40 ];
assign rho_out[1][2][ 20 ] = rho_in[1][2][ 14 ];
assign rho_out[1][3][ 20 ] = rho_in[1][3][ 29 ];
assign rho_out[1][4][ 20 ] = rho_in[1][4][ 0 ];
assign rho_out[2][0][ 20 ] = rho_in[2][0][ 17 ];
assign rho_out[2][1][ 20 ] = rho_in[2][1][ 10 ];
assign rho_out[2][2][ 20 ] = rho_in[2][2][ 41 ];
assign rho_out[2][3][ 20 ] = rho_in[2][3][ 59 ];
assign rho_out[2][4][ 20 ] = rho_in[2][4][ 45 ];
assign rho_out[3][0][ 20 ] = rho_in[3][0][ 43 ];
assign rho_out[3][1][ 20 ] = rho_in[3][1][ 39 ];
assign rho_out[3][2][ 20 ] = rho_in[3][2][ 5 ];
assign rho_out[3][3][ 20 ] = rho_in[3][3][ 63 ];
assign rho_out[3][4][ 20 ] = rho_in[3][4][ 12 ];
assign rho_out[4][0][ 20 ] = rho_in[4][0][ 2 ];
assign rho_out[4][1][ 20 ] = rho_in[4][1][ 18 ];
assign rho_out[4][2][ 20 ] = rho_in[4][2][ 23 ];
assign rho_out[4][3][ 20 ] = rho_in[4][3][ 28 ];
assign rho_out[4][4][ 20 ] = rho_in[4][4][ 6 ];
assign rho_out[0][0][ 21 ] = rho_in[0][0][ 21 ];
assign rho_out[0][1][ 21 ] = rho_in[0][1][ 20 ];
assign rho_out[0][2][ 21 ] = rho_in[0][2][ 23 ];
assign rho_out[0][3][ 21 ] = rho_in[0][3][ 57 ];
assign rho_out[0][4][ 21 ] = rho_in[0][4][ 58 ];
assign rho_out[1][0][ 21 ] = rho_in[1][0][ 49 ];
assign rho_out[1][1][ 21 ] = rho_in[1][1][ 41 ];
assign rho_out[1][2][ 21 ] = rho_in[1][2][ 15 ];
assign rho_out[1][3][ 21 ] = rho_in[1][3][ 30 ];
assign rho_out[1][4][ 21 ] = rho_in[1][4][ 1 ];
assign rho_out[2][0][ 21 ] = rho_in[2][0][ 18 ];
assign rho_out[2][1][ 21 ] = rho_in[2][1][ 11 ];
assign rho_out[2][2][ 21 ] = rho_in[2][2][ 42 ];
assign rho_out[2][3][ 21 ] = rho_in[2][3][ 60 ];
assign rho_out[2][4][ 21 ] = rho_in[2][4][ 46 ];
assign rho_out[3][0][ 21 ] = rho_in[3][0][ 44 ];
assign rho_out[3][1][ 21 ] = rho_in[3][1][ 40 ];
assign rho_out[3][2][ 21 ] = rho_in[3][2][ 6 ];
assign rho_out[3][3][ 21 ] = rho_in[3][3][ 0 ];
assign rho_out[3][4][ 21 ] = rho_in[3][4][ 13 ];
assign rho_out[4][0][ 21 ] = rho_in[4][0][ 3 ];
assign rho_out[4][1][ 21 ] = rho_in[4][1][ 19 ];
assign rho_out[4][2][ 21 ] = rho_in[4][2][ 24 ];
assign rho_out[4][3][ 21 ] = rho_in[4][3][ 29 ];
assign rho_out[4][4][ 21 ] = rho_in[4][4][ 7 ];
assign rho_out[0][0][ 22 ] = rho_in[0][0][ 22 ];
assign rho_out[0][1][ 22 ] = rho_in[0][1][ 21 ];
assign rho_out[0][2][ 22 ] = rho_in[0][2][ 24 ];
assign rho_out[0][3][ 22 ] = rho_in[0][3][ 58 ];
assign rho_out[0][4][ 22 ] = rho_in[0][4][ 59 ];
assign rho_out[1][0][ 22 ] = rho_in[1][0][ 50 ];
assign rho_out[1][1][ 22 ] = rho_in[1][1][ 42 ];
assign rho_out[1][2][ 22 ] = rho_in[1][2][ 16 ];
assign rho_out[1][3][ 22 ] = rho_in[1][3][ 31 ];
assign rho_out[1][4][ 22 ] = rho_in[1][4][ 2 ];
assign rho_out[2][0][ 22 ] = rho_in[2][0][ 19 ];
assign rho_out[2][1][ 22 ] = rho_in[2][1][ 12 ];
assign rho_out[2][2][ 22 ] = rho_in[2][2][ 43 ];
assign rho_out[2][3][ 22 ] = rho_in[2][3][ 61 ];
assign rho_out[2][4][ 22 ] = rho_in[2][4][ 47 ];
assign rho_out[3][0][ 22 ] = rho_in[3][0][ 45 ];
assign rho_out[3][1][ 22 ] = rho_in[3][1][ 41 ];
assign rho_out[3][2][ 22 ] = rho_in[3][2][ 7 ];
assign rho_out[3][3][ 22 ] = rho_in[3][3][ 1 ];
assign rho_out[3][4][ 22 ] = rho_in[3][4][ 14 ];
assign rho_out[4][0][ 22 ] = rho_in[4][0][ 4 ];
assign rho_out[4][1][ 22 ] = rho_in[4][1][ 20 ];
assign rho_out[4][2][ 22 ] = rho_in[4][2][ 25 ];
assign rho_out[4][3][ 22 ] = rho_in[4][3][ 30 ];
assign rho_out[4][4][ 22 ] = rho_in[4][4][ 8 ];
assign rho_out[0][0][ 23 ] = rho_in[0][0][ 23 ];
assign rho_out[0][1][ 23 ] = rho_in[0][1][ 22 ];
assign rho_out[0][2][ 23 ] = rho_in[0][2][ 25 ];
assign rho_out[0][3][ 23 ] = rho_in[0][3][ 59 ];
assign rho_out[0][4][ 23 ] = rho_in[0][4][ 60 ];
assign rho_out[1][0][ 23 ] = rho_in[1][0][ 51 ];
assign rho_out[1][1][ 23 ] = rho_in[1][1][ 43 ];
assign rho_out[1][2][ 23 ] = rho_in[1][2][ 17 ];
assign rho_out[1][3][ 23 ] = rho_in[1][3][ 32 ];
assign rho_out[1][4][ 23 ] = rho_in[1][4][ 3 ];
assign rho_out[2][0][ 23 ] = rho_in[2][0][ 20 ];
assign rho_out[2][1][ 23 ] = rho_in[2][1][ 13 ];
assign rho_out[2][2][ 23 ] = rho_in[2][2][ 44 ];
assign rho_out[2][3][ 23 ] = rho_in[2][3][ 62 ];
assign rho_out[2][4][ 23 ] = rho_in[2][4][ 48 ];
assign rho_out[3][0][ 23 ] = rho_in[3][0][ 46 ];
assign rho_out[3][1][ 23 ] = rho_in[3][1][ 42 ];
assign rho_out[3][2][ 23 ] = rho_in[3][2][ 8 ];
assign rho_out[3][3][ 23 ] = rho_in[3][3][ 2 ];
assign rho_out[3][4][ 23 ] = rho_in[3][4][ 15 ];
assign rho_out[4][0][ 23 ] = rho_in[4][0][ 5 ];
assign rho_out[4][1][ 23 ] = rho_in[4][1][ 21 ];
assign rho_out[4][2][ 23 ] = rho_in[4][2][ 26 ];
assign rho_out[4][3][ 23 ] = rho_in[4][3][ 31 ];
assign rho_out[4][4][ 23 ] = rho_in[4][4][ 9 ];
assign rho_out[0][0][ 24 ] = rho_in[0][0][ 24 ];
assign rho_out[0][1][ 24 ] = rho_in[0][1][ 23 ];
assign rho_out[0][2][ 24 ] = rho_in[0][2][ 26 ];
assign rho_out[0][3][ 24 ] = rho_in[0][3][ 60 ];
assign rho_out[0][4][ 24 ] = rho_in[0][4][ 61 ];
assign rho_out[1][0][ 24 ] = rho_in[1][0][ 52 ];
assign rho_out[1][1][ 24 ] = rho_in[1][1][ 44 ];
assign rho_out[1][2][ 24 ] = rho_in[1][2][ 18 ];
assign rho_out[1][3][ 24 ] = rho_in[1][3][ 33 ];
assign rho_out[1][4][ 24 ] = rho_in[1][4][ 4 ];
assign rho_out[2][0][ 24 ] = rho_in[2][0][ 21 ];
assign rho_out[2][1][ 24 ] = rho_in[2][1][ 14 ];
assign rho_out[2][2][ 24 ] = rho_in[2][2][ 45 ];
assign rho_out[2][3][ 24 ] = rho_in[2][3][ 63 ];
assign rho_out[2][4][ 24 ] = rho_in[2][4][ 49 ];
assign rho_out[3][0][ 24 ] = rho_in[3][0][ 47 ];
assign rho_out[3][1][ 24 ] = rho_in[3][1][ 43 ];
assign rho_out[3][2][ 24 ] = rho_in[3][2][ 9 ];
assign rho_out[3][3][ 24 ] = rho_in[3][3][ 3 ];
assign rho_out[3][4][ 24 ] = rho_in[3][4][ 16 ];
assign rho_out[4][0][ 24 ] = rho_in[4][0][ 6 ];
assign rho_out[4][1][ 24 ] = rho_in[4][1][ 22 ];
assign rho_out[4][2][ 24 ] = rho_in[4][2][ 27 ];
assign rho_out[4][3][ 24 ] = rho_in[4][3][ 32 ];
assign rho_out[4][4][ 24 ] = rho_in[4][4][ 10 ];
assign rho_out[0][0][ 25 ] = rho_in[0][0][ 25 ];
assign rho_out[0][1][ 25 ] = rho_in[0][1][ 24 ];
assign rho_out[0][2][ 25 ] = rho_in[0][2][ 27 ];
assign rho_out[0][3][ 25 ] = rho_in[0][3][ 61 ];
assign rho_out[0][4][ 25 ] = rho_in[0][4][ 62 ];
assign rho_out[1][0][ 25 ] = rho_in[1][0][ 53 ];
assign rho_out[1][1][ 25 ] = rho_in[1][1][ 45 ];
assign rho_out[1][2][ 25 ] = rho_in[1][2][ 19 ];
assign rho_out[1][3][ 25 ] = rho_in[1][3][ 34 ];
assign rho_out[1][4][ 25 ] = rho_in[1][4][ 5 ];
assign rho_out[2][0][ 25 ] = rho_in[2][0][ 22 ];
assign rho_out[2][1][ 25 ] = rho_in[2][1][ 15 ];
assign rho_out[2][2][ 25 ] = rho_in[2][2][ 46 ];
assign rho_out[2][3][ 25 ] = rho_in[2][3][ 0 ];
assign rho_out[2][4][ 25 ] = rho_in[2][4][ 50 ];
assign rho_out[3][0][ 25 ] = rho_in[3][0][ 48 ];
assign rho_out[3][1][ 25 ] = rho_in[3][1][ 44 ];
assign rho_out[3][2][ 25 ] = rho_in[3][2][ 10 ];
assign rho_out[3][3][ 25 ] = rho_in[3][3][ 4 ];
assign rho_out[3][4][ 25 ] = rho_in[3][4][ 17 ];
assign rho_out[4][0][ 25 ] = rho_in[4][0][ 7 ];
assign rho_out[4][1][ 25 ] = rho_in[4][1][ 23 ];
assign rho_out[4][2][ 25 ] = rho_in[4][2][ 28 ];
assign rho_out[4][3][ 25 ] = rho_in[4][3][ 33 ];
assign rho_out[4][4][ 25 ] = rho_in[4][4][ 11 ];
assign rho_out[0][0][ 26 ] = rho_in[0][0][ 26 ];
assign rho_out[0][1][ 26 ] = rho_in[0][1][ 25 ];
assign rho_out[0][2][ 26 ] = rho_in[0][2][ 28 ];
assign rho_out[0][3][ 26 ] = rho_in[0][3][ 62 ];
assign rho_out[0][4][ 26 ] = rho_in[0][4][ 63 ];
assign rho_out[1][0][ 26 ] = rho_in[1][0][ 54 ];
assign rho_out[1][1][ 26 ] = rho_in[1][1][ 46 ];
assign rho_out[1][2][ 26 ] = rho_in[1][2][ 20 ];
assign rho_out[1][3][ 26 ] = rho_in[1][3][ 35 ];
assign rho_out[1][4][ 26 ] = rho_in[1][4][ 6 ];
assign rho_out[2][0][ 26 ] = rho_in[2][0][ 23 ];
assign rho_out[2][1][ 26 ] = rho_in[2][1][ 16 ];
assign rho_out[2][2][ 26 ] = rho_in[2][2][ 47 ];
assign rho_out[2][3][ 26 ] = rho_in[2][3][ 1 ];
assign rho_out[2][4][ 26 ] = rho_in[2][4][ 51 ];
assign rho_out[3][0][ 26 ] = rho_in[3][0][ 49 ];
assign rho_out[3][1][ 26 ] = rho_in[3][1][ 45 ];
assign rho_out[3][2][ 26 ] = rho_in[3][2][ 11 ];
assign rho_out[3][3][ 26 ] = rho_in[3][3][ 5 ];
assign rho_out[3][4][ 26 ] = rho_in[3][4][ 18 ];
assign rho_out[4][0][ 26 ] = rho_in[4][0][ 8 ];
assign rho_out[4][1][ 26 ] = rho_in[4][1][ 24 ];
assign rho_out[4][2][ 26 ] = rho_in[4][2][ 29 ];
assign rho_out[4][3][ 26 ] = rho_in[4][3][ 34 ];
assign rho_out[4][4][ 26 ] = rho_in[4][4][ 12 ];
assign rho_out[0][0][ 27 ] = rho_in[0][0][ 27 ];
assign rho_out[0][1][ 27 ] = rho_in[0][1][ 26 ];
assign rho_out[0][2][ 27 ] = rho_in[0][2][ 29 ];
assign rho_out[0][3][ 27 ] = rho_in[0][3][ 63 ];
assign rho_out[0][4][ 27 ] = rho_in[0][4][ 0 ];
assign rho_out[1][0][ 27 ] = rho_in[1][0][ 55 ];
assign rho_out[1][1][ 27 ] = rho_in[1][1][ 47 ];
assign rho_out[1][2][ 27 ] = rho_in[1][2][ 21 ];
assign rho_out[1][3][ 27 ] = rho_in[1][3][ 36 ];
assign rho_out[1][4][ 27 ] = rho_in[1][4][ 7 ];
assign rho_out[2][0][ 27 ] = rho_in[2][0][ 24 ];
assign rho_out[2][1][ 27 ] = rho_in[2][1][ 17 ];
assign rho_out[2][2][ 27 ] = rho_in[2][2][ 48 ];
assign rho_out[2][3][ 27 ] = rho_in[2][3][ 2 ];
assign rho_out[2][4][ 27 ] = rho_in[2][4][ 52 ];
assign rho_out[3][0][ 27 ] = rho_in[3][0][ 50 ];
assign rho_out[3][1][ 27 ] = rho_in[3][1][ 46 ];
assign rho_out[3][2][ 27 ] = rho_in[3][2][ 12 ];
assign rho_out[3][3][ 27 ] = rho_in[3][3][ 6 ];
assign rho_out[3][4][ 27 ] = rho_in[3][4][ 19 ];
assign rho_out[4][0][ 27 ] = rho_in[4][0][ 9 ];
assign rho_out[4][1][ 27 ] = rho_in[4][1][ 25 ];
assign rho_out[4][2][ 27 ] = rho_in[4][2][ 30 ];
assign rho_out[4][3][ 27 ] = rho_in[4][3][ 35 ];
assign rho_out[4][4][ 27 ] = rho_in[4][4][ 13 ];
assign rho_out[0][0][ 28 ] = rho_in[0][0][ 28 ];
assign rho_out[0][1][ 28 ] = rho_in[0][1][ 27 ];
assign rho_out[0][2][ 28 ] = rho_in[0][2][ 30 ];
assign rho_out[0][3][ 28 ] = rho_in[0][3][ 0 ];
assign rho_out[0][4][ 28 ] = rho_in[0][4][ 1 ];
assign rho_out[1][0][ 28 ] = rho_in[1][0][ 56 ];
assign rho_out[1][1][ 28 ] = rho_in[1][1][ 48 ];
assign rho_out[1][2][ 28 ] = rho_in[1][2][ 22 ];
assign rho_out[1][3][ 28 ] = rho_in[1][3][ 37 ];
assign rho_out[1][4][ 28 ] = rho_in[1][4][ 8 ];
assign rho_out[2][0][ 28 ] = rho_in[2][0][ 25 ];
assign rho_out[2][1][ 28 ] = rho_in[2][1][ 18 ];
assign rho_out[2][2][ 28 ] = rho_in[2][2][ 49 ];
assign rho_out[2][3][ 28 ] = rho_in[2][3][ 3 ];
assign rho_out[2][4][ 28 ] = rho_in[2][4][ 53 ];
assign rho_out[3][0][ 28 ] = rho_in[3][0][ 51 ];
assign rho_out[3][1][ 28 ] = rho_in[3][1][ 47 ];
assign rho_out[3][2][ 28 ] = rho_in[3][2][ 13 ];
assign rho_out[3][3][ 28 ] = rho_in[3][3][ 7 ];
assign rho_out[3][4][ 28 ] = rho_in[3][4][ 20 ];
assign rho_out[4][0][ 28 ] = rho_in[4][0][ 10 ];
assign rho_out[4][1][ 28 ] = rho_in[4][1][ 26 ];
assign rho_out[4][2][ 28 ] = rho_in[4][2][ 31 ];
assign rho_out[4][3][ 28 ] = rho_in[4][3][ 36 ];
assign rho_out[4][4][ 28 ] = rho_in[4][4][ 14 ];
assign rho_out[0][0][ 29 ] = rho_in[0][0][ 29 ];
assign rho_out[0][1][ 29 ] = rho_in[0][1][ 28 ];
assign rho_out[0][2][ 29 ] = rho_in[0][2][ 31 ];
assign rho_out[0][3][ 29 ] = rho_in[0][3][ 1 ];
assign rho_out[0][4][ 29 ] = rho_in[0][4][ 2 ];
assign rho_out[1][0][ 29 ] = rho_in[1][0][ 57 ];
assign rho_out[1][1][ 29 ] = rho_in[1][1][ 49 ];
assign rho_out[1][2][ 29 ] = rho_in[1][2][ 23 ];
assign rho_out[1][3][ 29 ] = rho_in[1][3][ 38 ];
assign rho_out[1][4][ 29 ] = rho_in[1][4][ 9 ];
assign rho_out[2][0][ 29 ] = rho_in[2][0][ 26 ];
assign rho_out[2][1][ 29 ] = rho_in[2][1][ 19 ];
assign rho_out[2][2][ 29 ] = rho_in[2][2][ 50 ];
assign rho_out[2][3][ 29 ] = rho_in[2][3][ 4 ];
assign rho_out[2][4][ 29 ] = rho_in[2][4][ 54 ];
assign rho_out[3][0][ 29 ] = rho_in[3][0][ 52 ];
assign rho_out[3][1][ 29 ] = rho_in[3][1][ 48 ];
assign rho_out[3][2][ 29 ] = rho_in[3][2][ 14 ];
assign rho_out[3][3][ 29 ] = rho_in[3][3][ 8 ];
assign rho_out[3][4][ 29 ] = rho_in[3][4][ 21 ];
assign rho_out[4][0][ 29 ] = rho_in[4][0][ 11 ];
assign rho_out[4][1][ 29 ] = rho_in[4][1][ 27 ];
assign rho_out[4][2][ 29 ] = rho_in[4][2][ 32 ];
assign rho_out[4][3][ 29 ] = rho_in[4][3][ 37 ];
assign rho_out[4][4][ 29 ] = rho_in[4][4][ 15 ];
assign rho_out[0][0][ 30 ] = rho_in[0][0][ 30 ];
assign rho_out[0][1][ 30 ] = rho_in[0][1][ 29 ];
assign rho_out[0][2][ 30 ] = rho_in[0][2][ 32 ];
assign rho_out[0][3][ 30 ] = rho_in[0][3][ 2 ];
assign rho_out[0][4][ 30 ] = rho_in[0][4][ 3 ];
assign rho_out[1][0][ 30 ] = rho_in[1][0][ 58 ];
assign rho_out[1][1][ 30 ] = rho_in[1][1][ 50 ];
assign rho_out[1][2][ 30 ] = rho_in[1][2][ 24 ];
assign rho_out[1][3][ 30 ] = rho_in[1][3][ 39 ];
assign rho_out[1][4][ 30 ] = rho_in[1][4][ 10 ];
assign rho_out[2][0][ 30 ] = rho_in[2][0][ 27 ];
assign rho_out[2][1][ 30 ] = rho_in[2][1][ 20 ];
assign rho_out[2][2][ 30 ] = rho_in[2][2][ 51 ];
assign rho_out[2][3][ 30 ] = rho_in[2][3][ 5 ];
assign rho_out[2][4][ 30 ] = rho_in[2][4][ 55 ];
assign rho_out[3][0][ 30 ] = rho_in[3][0][ 53 ];
assign rho_out[3][1][ 30 ] = rho_in[3][1][ 49 ];
assign rho_out[3][2][ 30 ] = rho_in[3][2][ 15 ];
assign rho_out[3][3][ 30 ] = rho_in[3][3][ 9 ];
assign rho_out[3][4][ 30 ] = rho_in[3][4][ 22 ];
assign rho_out[4][0][ 30 ] = rho_in[4][0][ 12 ];
assign rho_out[4][1][ 30 ] = rho_in[4][1][ 28 ];
assign rho_out[4][2][ 30 ] = rho_in[4][2][ 33 ];
assign rho_out[4][3][ 30 ] = rho_in[4][3][ 38 ];
assign rho_out[4][4][ 30 ] = rho_in[4][4][ 16 ];
assign rho_out[0][0][ 31 ] = rho_in[0][0][ 31 ];
assign rho_out[0][1][ 31 ] = rho_in[0][1][ 30 ];
assign rho_out[0][2][ 31 ] = rho_in[0][2][ 33 ];
assign rho_out[0][3][ 31 ] = rho_in[0][3][ 3 ];
assign rho_out[0][4][ 31 ] = rho_in[0][4][ 4 ];
assign rho_out[1][0][ 31 ] = rho_in[1][0][ 59 ];
assign rho_out[1][1][ 31 ] = rho_in[1][1][ 51 ];
assign rho_out[1][2][ 31 ] = rho_in[1][2][ 25 ];
assign rho_out[1][3][ 31 ] = rho_in[1][3][ 40 ];
assign rho_out[1][4][ 31 ] = rho_in[1][4][ 11 ];
assign rho_out[2][0][ 31 ] = rho_in[2][0][ 28 ];
assign rho_out[2][1][ 31 ] = rho_in[2][1][ 21 ];
assign rho_out[2][2][ 31 ] = rho_in[2][2][ 52 ];
assign rho_out[2][3][ 31 ] = rho_in[2][3][ 6 ];
assign rho_out[2][4][ 31 ] = rho_in[2][4][ 56 ];
assign rho_out[3][0][ 31 ] = rho_in[3][0][ 54 ];
assign rho_out[3][1][ 31 ] = rho_in[3][1][ 50 ];
assign rho_out[3][2][ 31 ] = rho_in[3][2][ 16 ];
assign rho_out[3][3][ 31 ] = rho_in[3][3][ 10 ];
assign rho_out[3][4][ 31 ] = rho_in[3][4][ 23 ];
assign rho_out[4][0][ 31 ] = rho_in[4][0][ 13 ];
assign rho_out[4][1][ 31 ] = rho_in[4][1][ 29 ];
assign rho_out[4][2][ 31 ] = rho_in[4][2][ 34 ];
assign rho_out[4][3][ 31 ] = rho_in[4][3][ 39 ];
assign rho_out[4][4][ 31 ] = rho_in[4][4][ 17 ];
assign rho_out[0][0][ 32 ] = rho_in[0][0][ 32 ];
assign rho_out[0][1][ 32 ] = rho_in[0][1][ 31 ];
assign rho_out[0][2][ 32 ] = rho_in[0][2][ 34 ];
assign rho_out[0][3][ 32 ] = rho_in[0][3][ 4 ];
assign rho_out[0][4][ 32 ] = rho_in[0][4][ 5 ];
assign rho_out[1][0][ 32 ] = rho_in[1][0][ 60 ];
assign rho_out[1][1][ 32 ] = rho_in[1][1][ 52 ];
assign rho_out[1][2][ 32 ] = rho_in[1][2][ 26 ];
assign rho_out[1][3][ 32 ] = rho_in[1][3][ 41 ];
assign rho_out[1][4][ 32 ] = rho_in[1][4][ 12 ];
assign rho_out[2][0][ 32 ] = rho_in[2][0][ 29 ];
assign rho_out[2][1][ 32 ] = rho_in[2][1][ 22 ];
assign rho_out[2][2][ 32 ] = rho_in[2][2][ 53 ];
assign rho_out[2][3][ 32 ] = rho_in[2][3][ 7 ];
assign rho_out[2][4][ 32 ] = rho_in[2][4][ 57 ];
assign rho_out[3][0][ 32 ] = rho_in[3][0][ 55 ];
assign rho_out[3][1][ 32 ] = rho_in[3][1][ 51 ];
assign rho_out[3][2][ 32 ] = rho_in[3][2][ 17 ];
assign rho_out[3][3][ 32 ] = rho_in[3][3][ 11 ];
assign rho_out[3][4][ 32 ] = rho_in[3][4][ 24 ];
assign rho_out[4][0][ 32 ] = rho_in[4][0][ 14 ];
assign rho_out[4][1][ 32 ] = rho_in[4][1][ 30 ];
assign rho_out[4][2][ 32 ] = rho_in[4][2][ 35 ];
assign rho_out[4][3][ 32 ] = rho_in[4][3][ 40 ];
assign rho_out[4][4][ 32 ] = rho_in[4][4][ 18 ];
assign rho_out[0][0][ 33 ] = rho_in[0][0][ 33 ];
assign rho_out[0][1][ 33 ] = rho_in[0][1][ 32 ];
assign rho_out[0][2][ 33 ] = rho_in[0][2][ 35 ];
assign rho_out[0][3][ 33 ] = rho_in[0][3][ 5 ];
assign rho_out[0][4][ 33 ] = rho_in[0][4][ 6 ];
assign rho_out[1][0][ 33 ] = rho_in[1][0][ 61 ];
assign rho_out[1][1][ 33 ] = rho_in[1][1][ 53 ];
assign rho_out[1][2][ 33 ] = rho_in[1][2][ 27 ];
assign rho_out[1][3][ 33 ] = rho_in[1][3][ 42 ];
assign rho_out[1][4][ 33 ] = rho_in[1][4][ 13 ];
assign rho_out[2][0][ 33 ] = rho_in[2][0][ 30 ];
assign rho_out[2][1][ 33 ] = rho_in[2][1][ 23 ];
assign rho_out[2][2][ 33 ] = rho_in[2][2][ 54 ];
assign rho_out[2][3][ 33 ] = rho_in[2][3][ 8 ];
assign rho_out[2][4][ 33 ] = rho_in[2][4][ 58 ];
assign rho_out[3][0][ 33 ] = rho_in[3][0][ 56 ];
assign rho_out[3][1][ 33 ] = rho_in[3][1][ 52 ];
assign rho_out[3][2][ 33 ] = rho_in[3][2][ 18 ];
assign rho_out[3][3][ 33 ] = rho_in[3][3][ 12 ];
assign rho_out[3][4][ 33 ] = rho_in[3][4][ 25 ];
assign rho_out[4][0][ 33 ] = rho_in[4][0][ 15 ];
assign rho_out[4][1][ 33 ] = rho_in[4][1][ 31 ];
assign rho_out[4][2][ 33 ] = rho_in[4][2][ 36 ];
assign rho_out[4][3][ 33 ] = rho_in[4][3][ 41 ];
assign rho_out[4][4][ 33 ] = rho_in[4][4][ 19 ];
assign rho_out[0][0][ 34 ] = rho_in[0][0][ 34 ];
assign rho_out[0][1][ 34 ] = rho_in[0][1][ 33 ];
assign rho_out[0][2][ 34 ] = rho_in[0][2][ 36 ];
assign rho_out[0][3][ 34 ] = rho_in[0][3][ 6 ];
assign rho_out[0][4][ 34 ] = rho_in[0][4][ 7 ];
assign rho_out[1][0][ 34 ] = rho_in[1][0][ 62 ];
assign rho_out[1][1][ 34 ] = rho_in[1][1][ 54 ];
assign rho_out[1][2][ 34 ] = rho_in[1][2][ 28 ];
assign rho_out[1][3][ 34 ] = rho_in[1][3][ 43 ];
assign rho_out[1][4][ 34 ] = rho_in[1][4][ 14 ];
assign rho_out[2][0][ 34 ] = rho_in[2][0][ 31 ];
assign rho_out[2][1][ 34 ] = rho_in[2][1][ 24 ];
assign rho_out[2][2][ 34 ] = rho_in[2][2][ 55 ];
assign rho_out[2][3][ 34 ] = rho_in[2][3][ 9 ];
assign rho_out[2][4][ 34 ] = rho_in[2][4][ 59 ];
assign rho_out[3][0][ 34 ] = rho_in[3][0][ 57 ];
assign rho_out[3][1][ 34 ] = rho_in[3][1][ 53 ];
assign rho_out[3][2][ 34 ] = rho_in[3][2][ 19 ];
assign rho_out[3][3][ 34 ] = rho_in[3][3][ 13 ];
assign rho_out[3][4][ 34 ] = rho_in[3][4][ 26 ];
assign rho_out[4][0][ 34 ] = rho_in[4][0][ 16 ];
assign rho_out[4][1][ 34 ] = rho_in[4][1][ 32 ];
assign rho_out[4][2][ 34 ] = rho_in[4][2][ 37 ];
assign rho_out[4][3][ 34 ] = rho_in[4][3][ 42 ];
assign rho_out[4][4][ 34 ] = rho_in[4][4][ 20 ];
assign rho_out[0][0][ 35 ] = rho_in[0][0][ 35 ];
assign rho_out[0][1][ 35 ] = rho_in[0][1][ 34 ];
assign rho_out[0][2][ 35 ] = rho_in[0][2][ 37 ];
assign rho_out[0][3][ 35 ] = rho_in[0][3][ 7 ];
assign rho_out[0][4][ 35 ] = rho_in[0][4][ 8 ];
assign rho_out[1][0][ 35 ] = rho_in[1][0][ 63 ];
assign rho_out[1][1][ 35 ] = rho_in[1][1][ 55 ];
assign rho_out[1][2][ 35 ] = rho_in[1][2][ 29 ];
assign rho_out[1][3][ 35 ] = rho_in[1][3][ 44 ];
assign rho_out[1][4][ 35 ] = rho_in[1][4][ 15 ];
assign rho_out[2][0][ 35 ] = rho_in[2][0][ 32 ];
assign rho_out[2][1][ 35 ] = rho_in[2][1][ 25 ];
assign rho_out[2][2][ 35 ] = rho_in[2][2][ 56 ];
assign rho_out[2][3][ 35 ] = rho_in[2][3][ 10 ];
assign rho_out[2][4][ 35 ] = rho_in[2][4][ 60 ];
assign rho_out[3][0][ 35 ] = rho_in[3][0][ 58 ];
assign rho_out[3][1][ 35 ] = rho_in[3][1][ 54 ];
assign rho_out[3][2][ 35 ] = rho_in[3][2][ 20 ];
assign rho_out[3][3][ 35 ] = rho_in[3][3][ 14 ];
assign rho_out[3][4][ 35 ] = rho_in[3][4][ 27 ];
assign rho_out[4][0][ 35 ] = rho_in[4][0][ 17 ];
assign rho_out[4][1][ 35 ] = rho_in[4][1][ 33 ];
assign rho_out[4][2][ 35 ] = rho_in[4][2][ 38 ];
assign rho_out[4][3][ 35 ] = rho_in[4][3][ 43 ];
assign rho_out[4][4][ 35 ] = rho_in[4][4][ 21 ];
assign rho_out[0][0][ 36 ] = rho_in[0][0][ 36 ];
assign rho_out[0][1][ 36 ] = rho_in[0][1][ 35 ];
assign rho_out[0][2][ 36 ] = rho_in[0][2][ 38 ];
assign rho_out[0][3][ 36 ] = rho_in[0][3][ 8 ];
assign rho_out[0][4][ 36 ] = rho_in[0][4][ 9 ];
assign rho_out[1][0][ 36 ] = rho_in[1][0][ 0 ];
assign rho_out[1][1][ 36 ] = rho_in[1][1][ 56 ];
assign rho_out[1][2][ 36 ] = rho_in[1][2][ 30 ];
assign rho_out[1][3][ 36 ] = rho_in[1][3][ 45 ];
assign rho_out[1][4][ 36 ] = rho_in[1][4][ 16 ];
assign rho_out[2][0][ 36 ] = rho_in[2][0][ 33 ];
assign rho_out[2][1][ 36 ] = rho_in[2][1][ 26 ];
assign rho_out[2][2][ 36 ] = rho_in[2][2][ 57 ];
assign rho_out[2][3][ 36 ] = rho_in[2][3][ 11 ];
assign rho_out[2][4][ 36 ] = rho_in[2][4][ 61 ];
assign rho_out[3][0][ 36 ] = rho_in[3][0][ 59 ];
assign rho_out[3][1][ 36 ] = rho_in[3][1][ 55 ];
assign rho_out[3][2][ 36 ] = rho_in[3][2][ 21 ];
assign rho_out[3][3][ 36 ] = rho_in[3][3][ 15 ];
assign rho_out[3][4][ 36 ] = rho_in[3][4][ 28 ];
assign rho_out[4][0][ 36 ] = rho_in[4][0][ 18 ];
assign rho_out[4][1][ 36 ] = rho_in[4][1][ 34 ];
assign rho_out[4][2][ 36 ] = rho_in[4][2][ 39 ];
assign rho_out[4][3][ 36 ] = rho_in[4][3][ 44 ];
assign rho_out[4][4][ 36 ] = rho_in[4][4][ 22 ];
assign rho_out[0][0][ 37 ] = rho_in[0][0][ 37 ];
assign rho_out[0][1][ 37 ] = rho_in[0][1][ 36 ];
assign rho_out[0][2][ 37 ] = rho_in[0][2][ 39 ];
assign rho_out[0][3][ 37 ] = rho_in[0][3][ 9 ];
assign rho_out[0][4][ 37 ] = rho_in[0][4][ 10 ];
assign rho_out[1][0][ 37 ] = rho_in[1][0][ 1 ];
assign rho_out[1][1][ 37 ] = rho_in[1][1][ 57 ];
assign rho_out[1][2][ 37 ] = rho_in[1][2][ 31 ];
assign rho_out[1][3][ 37 ] = rho_in[1][3][ 46 ];
assign rho_out[1][4][ 37 ] = rho_in[1][4][ 17 ];
assign rho_out[2][0][ 37 ] = rho_in[2][0][ 34 ];
assign rho_out[2][1][ 37 ] = rho_in[2][1][ 27 ];
assign rho_out[2][2][ 37 ] = rho_in[2][2][ 58 ];
assign rho_out[2][3][ 37 ] = rho_in[2][3][ 12 ];
assign rho_out[2][4][ 37 ] = rho_in[2][4][ 62 ];
assign rho_out[3][0][ 37 ] = rho_in[3][0][ 60 ];
assign rho_out[3][1][ 37 ] = rho_in[3][1][ 56 ];
assign rho_out[3][2][ 37 ] = rho_in[3][2][ 22 ];
assign rho_out[3][3][ 37 ] = rho_in[3][3][ 16 ];
assign rho_out[3][4][ 37 ] = rho_in[3][4][ 29 ];
assign rho_out[4][0][ 37 ] = rho_in[4][0][ 19 ];
assign rho_out[4][1][ 37 ] = rho_in[4][1][ 35 ];
assign rho_out[4][2][ 37 ] = rho_in[4][2][ 40 ];
assign rho_out[4][3][ 37 ] = rho_in[4][3][ 45 ];
assign rho_out[4][4][ 37 ] = rho_in[4][4][ 23 ];
assign rho_out[0][0][ 38 ] = rho_in[0][0][ 38 ];
assign rho_out[0][1][ 38 ] = rho_in[0][1][ 37 ];
assign rho_out[0][2][ 38 ] = rho_in[0][2][ 40 ];
assign rho_out[0][3][ 38 ] = rho_in[0][3][ 10 ];
assign rho_out[0][4][ 38 ] = rho_in[0][4][ 11 ];
assign rho_out[1][0][ 38 ] = rho_in[1][0][ 2 ];
assign rho_out[1][1][ 38 ] = rho_in[1][1][ 58 ];
assign rho_out[1][2][ 38 ] = rho_in[1][2][ 32 ];
assign rho_out[1][3][ 38 ] = rho_in[1][3][ 47 ];
assign rho_out[1][4][ 38 ] = rho_in[1][4][ 18 ];
assign rho_out[2][0][ 38 ] = rho_in[2][0][ 35 ];
assign rho_out[2][1][ 38 ] = rho_in[2][1][ 28 ];
assign rho_out[2][2][ 38 ] = rho_in[2][2][ 59 ];
assign rho_out[2][3][ 38 ] = rho_in[2][3][ 13 ];
assign rho_out[2][4][ 38 ] = rho_in[2][4][ 63 ];
assign rho_out[3][0][ 38 ] = rho_in[3][0][ 61 ];
assign rho_out[3][1][ 38 ] = rho_in[3][1][ 57 ];
assign rho_out[3][2][ 38 ] = rho_in[3][2][ 23 ];
assign rho_out[3][3][ 38 ] = rho_in[3][3][ 17 ];
assign rho_out[3][4][ 38 ] = rho_in[3][4][ 30 ];
assign rho_out[4][0][ 38 ] = rho_in[4][0][ 20 ];
assign rho_out[4][1][ 38 ] = rho_in[4][1][ 36 ];
assign rho_out[4][2][ 38 ] = rho_in[4][2][ 41 ];
assign rho_out[4][3][ 38 ] = rho_in[4][3][ 46 ];
assign rho_out[4][4][ 38 ] = rho_in[4][4][ 24 ];
assign rho_out[0][0][ 39 ] = rho_in[0][0][ 39 ];
assign rho_out[0][1][ 39 ] = rho_in[0][1][ 38 ];
assign rho_out[0][2][ 39 ] = rho_in[0][2][ 41 ];
assign rho_out[0][3][ 39 ] = rho_in[0][3][ 11 ];
assign rho_out[0][4][ 39 ] = rho_in[0][4][ 12 ];
assign rho_out[1][0][ 39 ] = rho_in[1][0][ 3 ];
assign rho_out[1][1][ 39 ] = rho_in[1][1][ 59 ];
assign rho_out[1][2][ 39 ] = rho_in[1][2][ 33 ];
assign rho_out[1][3][ 39 ] = rho_in[1][3][ 48 ];
assign rho_out[1][4][ 39 ] = rho_in[1][4][ 19 ];
assign rho_out[2][0][ 39 ] = rho_in[2][0][ 36 ];
assign rho_out[2][1][ 39 ] = rho_in[2][1][ 29 ];
assign rho_out[2][2][ 39 ] = rho_in[2][2][ 60 ];
assign rho_out[2][3][ 39 ] = rho_in[2][3][ 14 ];
assign rho_out[2][4][ 39 ] = rho_in[2][4][ 0 ];
assign rho_out[3][0][ 39 ] = rho_in[3][0][ 62 ];
assign rho_out[3][1][ 39 ] = rho_in[3][1][ 58 ];
assign rho_out[3][2][ 39 ] = rho_in[3][2][ 24 ];
assign rho_out[3][3][ 39 ] = rho_in[3][3][ 18 ];
assign rho_out[3][4][ 39 ] = rho_in[3][4][ 31 ];
assign rho_out[4][0][ 39 ] = rho_in[4][0][ 21 ];
assign rho_out[4][1][ 39 ] = rho_in[4][1][ 37 ];
assign rho_out[4][2][ 39 ] = rho_in[4][2][ 42 ];
assign rho_out[4][3][ 39 ] = rho_in[4][3][ 47 ];
assign rho_out[4][4][ 39 ] = rho_in[4][4][ 25 ];
assign rho_out[0][0][ 40 ] = rho_in[0][0][ 40 ];
assign rho_out[0][1][ 40 ] = rho_in[0][1][ 39 ];
assign rho_out[0][2][ 40 ] = rho_in[0][2][ 42 ];
assign rho_out[0][3][ 40 ] = rho_in[0][3][ 12 ];
assign rho_out[0][4][ 40 ] = rho_in[0][4][ 13 ];
assign rho_out[1][0][ 40 ] = rho_in[1][0][ 4 ];
assign rho_out[1][1][ 40 ] = rho_in[1][1][ 60 ];
assign rho_out[1][2][ 40 ] = rho_in[1][2][ 34 ];
assign rho_out[1][3][ 40 ] = rho_in[1][3][ 49 ];
assign rho_out[1][4][ 40 ] = rho_in[1][4][ 20 ];
assign rho_out[2][0][ 40 ] = rho_in[2][0][ 37 ];
assign rho_out[2][1][ 40 ] = rho_in[2][1][ 30 ];
assign rho_out[2][2][ 40 ] = rho_in[2][2][ 61 ];
assign rho_out[2][3][ 40 ] = rho_in[2][3][ 15 ];
assign rho_out[2][4][ 40 ] = rho_in[2][4][ 1 ];
assign rho_out[3][0][ 40 ] = rho_in[3][0][ 63 ];
assign rho_out[3][1][ 40 ] = rho_in[3][1][ 59 ];
assign rho_out[3][2][ 40 ] = rho_in[3][2][ 25 ];
assign rho_out[3][3][ 40 ] = rho_in[3][3][ 19 ];
assign rho_out[3][4][ 40 ] = rho_in[3][4][ 32 ];
assign rho_out[4][0][ 40 ] = rho_in[4][0][ 22 ];
assign rho_out[4][1][ 40 ] = rho_in[4][1][ 38 ];
assign rho_out[4][2][ 40 ] = rho_in[4][2][ 43 ];
assign rho_out[4][3][ 40 ] = rho_in[4][3][ 48 ];
assign rho_out[4][4][ 40 ] = rho_in[4][4][ 26 ];
assign rho_out[0][0][ 41 ] = rho_in[0][0][ 41 ];
assign rho_out[0][1][ 41 ] = rho_in[0][1][ 40 ];
assign rho_out[0][2][ 41 ] = rho_in[0][2][ 43 ];
assign rho_out[0][3][ 41 ] = rho_in[0][3][ 13 ];
assign rho_out[0][4][ 41 ] = rho_in[0][4][ 14 ];
assign rho_out[1][0][ 41 ] = rho_in[1][0][ 5 ];
assign rho_out[1][1][ 41 ] = rho_in[1][1][ 61 ];
assign rho_out[1][2][ 41 ] = rho_in[1][2][ 35 ];
assign rho_out[1][3][ 41 ] = rho_in[1][3][ 50 ];
assign rho_out[1][4][ 41 ] = rho_in[1][4][ 21 ];
assign rho_out[2][0][ 41 ] = rho_in[2][0][ 38 ];
assign rho_out[2][1][ 41 ] = rho_in[2][1][ 31 ];
assign rho_out[2][2][ 41 ] = rho_in[2][2][ 62 ];
assign rho_out[2][3][ 41 ] = rho_in[2][3][ 16 ];
assign rho_out[2][4][ 41 ] = rho_in[2][4][ 2 ];
assign rho_out[3][0][ 41 ] = rho_in[3][0][ 0 ];
assign rho_out[3][1][ 41 ] = rho_in[3][1][ 60 ];
assign rho_out[3][2][ 41 ] = rho_in[3][2][ 26 ];
assign rho_out[3][3][ 41 ] = rho_in[3][3][ 20 ];
assign rho_out[3][4][ 41 ] = rho_in[3][4][ 33 ];
assign rho_out[4][0][ 41 ] = rho_in[4][0][ 23 ];
assign rho_out[4][1][ 41 ] = rho_in[4][1][ 39 ];
assign rho_out[4][2][ 41 ] = rho_in[4][2][ 44 ];
assign rho_out[4][3][ 41 ] = rho_in[4][3][ 49 ];
assign rho_out[4][4][ 41 ] = rho_in[4][4][ 27 ];
assign rho_out[0][0][ 42 ] = rho_in[0][0][ 42 ];
assign rho_out[0][1][ 42 ] = rho_in[0][1][ 41 ];
assign rho_out[0][2][ 42 ] = rho_in[0][2][ 44 ];
assign rho_out[0][3][ 42 ] = rho_in[0][3][ 14 ];
assign rho_out[0][4][ 42 ] = rho_in[0][4][ 15 ];
assign rho_out[1][0][ 42 ] = rho_in[1][0][ 6 ];
assign rho_out[1][1][ 42 ] = rho_in[1][1][ 62 ];
assign rho_out[1][2][ 42 ] = rho_in[1][2][ 36 ];
assign rho_out[1][3][ 42 ] = rho_in[1][3][ 51 ];
assign rho_out[1][4][ 42 ] = rho_in[1][4][ 22 ];
assign rho_out[2][0][ 42 ] = rho_in[2][0][ 39 ];
assign rho_out[2][1][ 42 ] = rho_in[2][1][ 32 ];
assign rho_out[2][2][ 42 ] = rho_in[2][2][ 63 ];
assign rho_out[2][3][ 42 ] = rho_in[2][3][ 17 ];
assign rho_out[2][4][ 42 ] = rho_in[2][4][ 3 ];
assign rho_out[3][0][ 42 ] = rho_in[3][0][ 1 ];
assign rho_out[3][1][ 42 ] = rho_in[3][1][ 61 ];
assign rho_out[3][2][ 42 ] = rho_in[3][2][ 27 ];
assign rho_out[3][3][ 42 ] = rho_in[3][3][ 21 ];
assign rho_out[3][4][ 42 ] = rho_in[3][4][ 34 ];
assign rho_out[4][0][ 42 ] = rho_in[4][0][ 24 ];
assign rho_out[4][1][ 42 ] = rho_in[4][1][ 40 ];
assign rho_out[4][2][ 42 ] = rho_in[4][2][ 45 ];
assign rho_out[4][3][ 42 ] = rho_in[4][3][ 50 ];
assign rho_out[4][4][ 42 ] = rho_in[4][4][ 28 ];
assign rho_out[0][0][ 43 ] = rho_in[0][0][ 43 ];
assign rho_out[0][1][ 43 ] = rho_in[0][1][ 42 ];
assign rho_out[0][2][ 43 ] = rho_in[0][2][ 45 ];
assign rho_out[0][3][ 43 ] = rho_in[0][3][ 15 ];
assign rho_out[0][4][ 43 ] = rho_in[0][4][ 16 ];
assign rho_out[1][0][ 43 ] = rho_in[1][0][ 7 ];
assign rho_out[1][1][ 43 ] = rho_in[1][1][ 63 ];
assign rho_out[1][2][ 43 ] = rho_in[1][2][ 37 ];
assign rho_out[1][3][ 43 ] = rho_in[1][3][ 52 ];
assign rho_out[1][4][ 43 ] = rho_in[1][4][ 23 ];
assign rho_out[2][0][ 43 ] = rho_in[2][0][ 40 ];
assign rho_out[2][1][ 43 ] = rho_in[2][1][ 33 ];
assign rho_out[2][2][ 43 ] = rho_in[2][2][ 0 ];
assign rho_out[2][3][ 43 ] = rho_in[2][3][ 18 ];
assign rho_out[2][4][ 43 ] = rho_in[2][4][ 4 ];
assign rho_out[3][0][ 43 ] = rho_in[3][0][ 2 ];
assign rho_out[3][1][ 43 ] = rho_in[3][1][ 62 ];
assign rho_out[3][2][ 43 ] = rho_in[3][2][ 28 ];
assign rho_out[3][3][ 43 ] = rho_in[3][3][ 22 ];
assign rho_out[3][4][ 43 ] = rho_in[3][4][ 35 ];
assign rho_out[4][0][ 43 ] = rho_in[4][0][ 25 ];
assign rho_out[4][1][ 43 ] = rho_in[4][1][ 41 ];
assign rho_out[4][2][ 43 ] = rho_in[4][2][ 46 ];
assign rho_out[4][3][ 43 ] = rho_in[4][3][ 51 ];
assign rho_out[4][4][ 43 ] = rho_in[4][4][ 29 ];
assign rho_out[0][0][ 44 ] = rho_in[0][0][ 44 ];
assign rho_out[0][1][ 44 ] = rho_in[0][1][ 43 ];
assign rho_out[0][2][ 44 ] = rho_in[0][2][ 46 ];
assign rho_out[0][3][ 44 ] = rho_in[0][3][ 16 ];
assign rho_out[0][4][ 44 ] = rho_in[0][4][ 17 ];
assign rho_out[1][0][ 44 ] = rho_in[1][0][ 8 ];
assign rho_out[1][1][ 44 ] = rho_in[1][1][ 0 ];
assign rho_out[1][2][ 44 ] = rho_in[1][2][ 38 ];
assign rho_out[1][3][ 44 ] = rho_in[1][3][ 53 ];
assign rho_out[1][4][ 44 ] = rho_in[1][4][ 24 ];
assign rho_out[2][0][ 44 ] = rho_in[2][0][ 41 ];
assign rho_out[2][1][ 44 ] = rho_in[2][1][ 34 ];
assign rho_out[2][2][ 44 ] = rho_in[2][2][ 1 ];
assign rho_out[2][3][ 44 ] = rho_in[2][3][ 19 ];
assign rho_out[2][4][ 44 ] = rho_in[2][4][ 5 ];
assign rho_out[3][0][ 44 ] = rho_in[3][0][ 3 ];
assign rho_out[3][1][ 44 ] = rho_in[3][1][ 63 ];
assign rho_out[3][2][ 44 ] = rho_in[3][2][ 29 ];
assign rho_out[3][3][ 44 ] = rho_in[3][3][ 23 ];
assign rho_out[3][4][ 44 ] = rho_in[3][4][ 36 ];
assign rho_out[4][0][ 44 ] = rho_in[4][0][ 26 ];
assign rho_out[4][1][ 44 ] = rho_in[4][1][ 42 ];
assign rho_out[4][2][ 44 ] = rho_in[4][2][ 47 ];
assign rho_out[4][3][ 44 ] = rho_in[4][3][ 52 ];
assign rho_out[4][4][ 44 ] = rho_in[4][4][ 30 ];
assign rho_out[0][0][ 45 ] = rho_in[0][0][ 45 ];
assign rho_out[0][1][ 45 ] = rho_in[0][1][ 44 ];
assign rho_out[0][2][ 45 ] = rho_in[0][2][ 47 ];
assign rho_out[0][3][ 45 ] = rho_in[0][3][ 17 ];
assign rho_out[0][4][ 45 ] = rho_in[0][4][ 18 ];
assign rho_out[1][0][ 45 ] = rho_in[1][0][ 9 ];
assign rho_out[1][1][ 45 ] = rho_in[1][1][ 1 ];
assign rho_out[1][2][ 45 ] = rho_in[1][2][ 39 ];
assign rho_out[1][3][ 45 ] = rho_in[1][3][ 54 ];
assign rho_out[1][4][ 45 ] = rho_in[1][4][ 25 ];
assign rho_out[2][0][ 45 ] = rho_in[2][0][ 42 ];
assign rho_out[2][1][ 45 ] = rho_in[2][1][ 35 ];
assign rho_out[2][2][ 45 ] = rho_in[2][2][ 2 ];
assign rho_out[2][3][ 45 ] = rho_in[2][3][ 20 ];
assign rho_out[2][4][ 45 ] = rho_in[2][4][ 6 ];
assign rho_out[3][0][ 45 ] = rho_in[3][0][ 4 ];
assign rho_out[3][1][ 45 ] = rho_in[3][1][ 0 ];
assign rho_out[3][2][ 45 ] = rho_in[3][2][ 30 ];
assign rho_out[3][3][ 45 ] = rho_in[3][3][ 24 ];
assign rho_out[3][4][ 45 ] = rho_in[3][4][ 37 ];
assign rho_out[4][0][ 45 ] = rho_in[4][0][ 27 ];
assign rho_out[4][1][ 45 ] = rho_in[4][1][ 43 ];
assign rho_out[4][2][ 45 ] = rho_in[4][2][ 48 ];
assign rho_out[4][3][ 45 ] = rho_in[4][3][ 53 ];
assign rho_out[4][4][ 45 ] = rho_in[4][4][ 31 ];
assign rho_out[0][0][ 46 ] = rho_in[0][0][ 46 ];
assign rho_out[0][1][ 46 ] = rho_in[0][1][ 45 ];
assign rho_out[0][2][ 46 ] = rho_in[0][2][ 48 ];
assign rho_out[0][3][ 46 ] = rho_in[0][3][ 18 ];
assign rho_out[0][4][ 46 ] = rho_in[0][4][ 19 ];
assign rho_out[1][0][ 46 ] = rho_in[1][0][ 10 ];
assign rho_out[1][1][ 46 ] = rho_in[1][1][ 2 ];
assign rho_out[1][2][ 46 ] = rho_in[1][2][ 40 ];
assign rho_out[1][3][ 46 ] = rho_in[1][3][ 55 ];
assign rho_out[1][4][ 46 ] = rho_in[1][4][ 26 ];
assign rho_out[2][0][ 46 ] = rho_in[2][0][ 43 ];
assign rho_out[2][1][ 46 ] = rho_in[2][1][ 36 ];
assign rho_out[2][2][ 46 ] = rho_in[2][2][ 3 ];
assign rho_out[2][3][ 46 ] = rho_in[2][3][ 21 ];
assign rho_out[2][4][ 46 ] = rho_in[2][4][ 7 ];
assign rho_out[3][0][ 46 ] = rho_in[3][0][ 5 ];
assign rho_out[3][1][ 46 ] = rho_in[3][1][ 1 ];
assign rho_out[3][2][ 46 ] = rho_in[3][2][ 31 ];
assign rho_out[3][3][ 46 ] = rho_in[3][3][ 25 ];
assign rho_out[3][4][ 46 ] = rho_in[3][4][ 38 ];
assign rho_out[4][0][ 46 ] = rho_in[4][0][ 28 ];
assign rho_out[4][1][ 46 ] = rho_in[4][1][ 44 ];
assign rho_out[4][2][ 46 ] = rho_in[4][2][ 49 ];
assign rho_out[4][3][ 46 ] = rho_in[4][3][ 54 ];
assign rho_out[4][4][ 46 ] = rho_in[4][4][ 32 ];
assign rho_out[0][0][ 47 ] = rho_in[0][0][ 47 ];
assign rho_out[0][1][ 47 ] = rho_in[0][1][ 46 ];
assign rho_out[0][2][ 47 ] = rho_in[0][2][ 49 ];
assign rho_out[0][3][ 47 ] = rho_in[0][3][ 19 ];
assign rho_out[0][4][ 47 ] = rho_in[0][4][ 20 ];
assign rho_out[1][0][ 47 ] = rho_in[1][0][ 11 ];
assign rho_out[1][1][ 47 ] = rho_in[1][1][ 3 ];
assign rho_out[1][2][ 47 ] = rho_in[1][2][ 41 ];
assign rho_out[1][3][ 47 ] = rho_in[1][3][ 56 ];
assign rho_out[1][4][ 47 ] = rho_in[1][4][ 27 ];
assign rho_out[2][0][ 47 ] = rho_in[2][0][ 44 ];
assign rho_out[2][1][ 47 ] = rho_in[2][1][ 37 ];
assign rho_out[2][2][ 47 ] = rho_in[2][2][ 4 ];
assign rho_out[2][3][ 47 ] = rho_in[2][3][ 22 ];
assign rho_out[2][4][ 47 ] = rho_in[2][4][ 8 ];
assign rho_out[3][0][ 47 ] = rho_in[3][0][ 6 ];
assign rho_out[3][1][ 47 ] = rho_in[3][1][ 2 ];
assign rho_out[3][2][ 47 ] = rho_in[3][2][ 32 ];
assign rho_out[3][3][ 47 ] = rho_in[3][3][ 26 ];
assign rho_out[3][4][ 47 ] = rho_in[3][4][ 39 ];
assign rho_out[4][0][ 47 ] = rho_in[4][0][ 29 ];
assign rho_out[4][1][ 47 ] = rho_in[4][1][ 45 ];
assign rho_out[4][2][ 47 ] = rho_in[4][2][ 50 ];
assign rho_out[4][3][ 47 ] = rho_in[4][3][ 55 ];
assign rho_out[4][4][ 47 ] = rho_in[4][4][ 33 ];
assign rho_out[0][0][ 48 ] = rho_in[0][0][ 48 ];
assign rho_out[0][1][ 48 ] = rho_in[0][1][ 47 ];
assign rho_out[0][2][ 48 ] = rho_in[0][2][ 50 ];
assign rho_out[0][3][ 48 ] = rho_in[0][3][ 20 ];
assign rho_out[0][4][ 48 ] = rho_in[0][4][ 21 ];
assign rho_out[1][0][ 48 ] = rho_in[1][0][ 12 ];
assign rho_out[1][1][ 48 ] = rho_in[1][1][ 4 ];
assign rho_out[1][2][ 48 ] = rho_in[1][2][ 42 ];
assign rho_out[1][3][ 48 ] = rho_in[1][3][ 57 ];
assign rho_out[1][4][ 48 ] = rho_in[1][4][ 28 ];
assign rho_out[2][0][ 48 ] = rho_in[2][0][ 45 ];
assign rho_out[2][1][ 48 ] = rho_in[2][1][ 38 ];
assign rho_out[2][2][ 48 ] = rho_in[2][2][ 5 ];
assign rho_out[2][3][ 48 ] = rho_in[2][3][ 23 ];
assign rho_out[2][4][ 48 ] = rho_in[2][4][ 9 ];
assign rho_out[3][0][ 48 ] = rho_in[3][0][ 7 ];
assign rho_out[3][1][ 48 ] = rho_in[3][1][ 3 ];
assign rho_out[3][2][ 48 ] = rho_in[3][2][ 33 ];
assign rho_out[3][3][ 48 ] = rho_in[3][3][ 27 ];
assign rho_out[3][4][ 48 ] = rho_in[3][4][ 40 ];
assign rho_out[4][0][ 48 ] = rho_in[4][0][ 30 ];
assign rho_out[4][1][ 48 ] = rho_in[4][1][ 46 ];
assign rho_out[4][2][ 48 ] = rho_in[4][2][ 51 ];
assign rho_out[4][3][ 48 ] = rho_in[4][3][ 56 ];
assign rho_out[4][4][ 48 ] = rho_in[4][4][ 34 ];
assign rho_out[0][0][ 49 ] = rho_in[0][0][ 49 ];
assign rho_out[0][1][ 49 ] = rho_in[0][1][ 48 ];
assign rho_out[0][2][ 49 ] = rho_in[0][2][ 51 ];
assign rho_out[0][3][ 49 ] = rho_in[0][3][ 21 ];
assign rho_out[0][4][ 49 ] = rho_in[0][4][ 22 ];
assign rho_out[1][0][ 49 ] = rho_in[1][0][ 13 ];
assign rho_out[1][1][ 49 ] = rho_in[1][1][ 5 ];
assign rho_out[1][2][ 49 ] = rho_in[1][2][ 43 ];
assign rho_out[1][3][ 49 ] = rho_in[1][3][ 58 ];
assign rho_out[1][4][ 49 ] = rho_in[1][4][ 29 ];
assign rho_out[2][0][ 49 ] = rho_in[2][0][ 46 ];
assign rho_out[2][1][ 49 ] = rho_in[2][1][ 39 ];
assign rho_out[2][2][ 49 ] = rho_in[2][2][ 6 ];
assign rho_out[2][3][ 49 ] = rho_in[2][3][ 24 ];
assign rho_out[2][4][ 49 ] = rho_in[2][4][ 10 ];
assign rho_out[3][0][ 49 ] = rho_in[3][0][ 8 ];
assign rho_out[3][1][ 49 ] = rho_in[3][1][ 4 ];
assign rho_out[3][2][ 49 ] = rho_in[3][2][ 34 ];
assign rho_out[3][3][ 49 ] = rho_in[3][3][ 28 ];
assign rho_out[3][4][ 49 ] = rho_in[3][4][ 41 ];
assign rho_out[4][0][ 49 ] = rho_in[4][0][ 31 ];
assign rho_out[4][1][ 49 ] = rho_in[4][1][ 47 ];
assign rho_out[4][2][ 49 ] = rho_in[4][2][ 52 ];
assign rho_out[4][3][ 49 ] = rho_in[4][3][ 57 ];
assign rho_out[4][4][ 49 ] = rho_in[4][4][ 35 ];
assign rho_out[0][0][ 50 ] = rho_in[0][0][ 50 ];
assign rho_out[0][1][ 50 ] = rho_in[0][1][ 49 ];
assign rho_out[0][2][ 50 ] = rho_in[0][2][ 52 ];
assign rho_out[0][3][ 50 ] = rho_in[0][3][ 22 ];
assign rho_out[0][4][ 50 ] = rho_in[0][4][ 23 ];
assign rho_out[1][0][ 50 ] = rho_in[1][0][ 14 ];
assign rho_out[1][1][ 50 ] = rho_in[1][1][ 6 ];
assign rho_out[1][2][ 50 ] = rho_in[1][2][ 44 ];
assign rho_out[1][3][ 50 ] = rho_in[1][3][ 59 ];
assign rho_out[1][4][ 50 ] = rho_in[1][4][ 30 ];
assign rho_out[2][0][ 50 ] = rho_in[2][0][ 47 ];
assign rho_out[2][1][ 50 ] = rho_in[2][1][ 40 ];
assign rho_out[2][2][ 50 ] = rho_in[2][2][ 7 ];
assign rho_out[2][3][ 50 ] = rho_in[2][3][ 25 ];
assign rho_out[2][4][ 50 ] = rho_in[2][4][ 11 ];
assign rho_out[3][0][ 50 ] = rho_in[3][0][ 9 ];
assign rho_out[3][1][ 50 ] = rho_in[3][1][ 5 ];
assign rho_out[3][2][ 50 ] = rho_in[3][2][ 35 ];
assign rho_out[3][3][ 50 ] = rho_in[3][3][ 29 ];
assign rho_out[3][4][ 50 ] = rho_in[3][4][ 42 ];
assign rho_out[4][0][ 50 ] = rho_in[4][0][ 32 ];
assign rho_out[4][1][ 50 ] = rho_in[4][1][ 48 ];
assign rho_out[4][2][ 50 ] = rho_in[4][2][ 53 ];
assign rho_out[4][3][ 50 ] = rho_in[4][3][ 58 ];
assign rho_out[4][4][ 50 ] = rho_in[4][4][ 36 ];
assign rho_out[0][0][ 51 ] = rho_in[0][0][ 51 ];
assign rho_out[0][1][ 51 ] = rho_in[0][1][ 50 ];
assign rho_out[0][2][ 51 ] = rho_in[0][2][ 53 ];
assign rho_out[0][3][ 51 ] = rho_in[0][3][ 23 ];
assign rho_out[0][4][ 51 ] = rho_in[0][4][ 24 ];
assign rho_out[1][0][ 51 ] = rho_in[1][0][ 15 ];
assign rho_out[1][1][ 51 ] = rho_in[1][1][ 7 ];
assign rho_out[1][2][ 51 ] = rho_in[1][2][ 45 ];
assign rho_out[1][3][ 51 ] = rho_in[1][3][ 60 ];
assign rho_out[1][4][ 51 ] = rho_in[1][4][ 31 ];
assign rho_out[2][0][ 51 ] = rho_in[2][0][ 48 ];
assign rho_out[2][1][ 51 ] = rho_in[2][1][ 41 ];
assign rho_out[2][2][ 51 ] = rho_in[2][2][ 8 ];
assign rho_out[2][3][ 51 ] = rho_in[2][3][ 26 ];
assign rho_out[2][4][ 51 ] = rho_in[2][4][ 12 ];
assign rho_out[3][0][ 51 ] = rho_in[3][0][ 10 ];
assign rho_out[3][1][ 51 ] = rho_in[3][1][ 6 ];
assign rho_out[3][2][ 51 ] = rho_in[3][2][ 36 ];
assign rho_out[3][3][ 51 ] = rho_in[3][3][ 30 ];
assign rho_out[3][4][ 51 ] = rho_in[3][4][ 43 ];
assign rho_out[4][0][ 51 ] = rho_in[4][0][ 33 ];
assign rho_out[4][1][ 51 ] = rho_in[4][1][ 49 ];
assign rho_out[4][2][ 51 ] = rho_in[4][2][ 54 ];
assign rho_out[4][3][ 51 ] = rho_in[4][3][ 59 ];
assign rho_out[4][4][ 51 ] = rho_in[4][4][ 37 ];
assign rho_out[0][0][ 52 ] = rho_in[0][0][ 52 ];
assign rho_out[0][1][ 52 ] = rho_in[0][1][ 51 ];
assign rho_out[0][2][ 52 ] = rho_in[0][2][ 54 ];
assign rho_out[0][3][ 52 ] = rho_in[0][3][ 24 ];
assign rho_out[0][4][ 52 ] = rho_in[0][4][ 25 ];
assign rho_out[1][0][ 52 ] = rho_in[1][0][ 16 ];
assign rho_out[1][1][ 52 ] = rho_in[1][1][ 8 ];
assign rho_out[1][2][ 52 ] = rho_in[1][2][ 46 ];
assign rho_out[1][3][ 52 ] = rho_in[1][3][ 61 ];
assign rho_out[1][4][ 52 ] = rho_in[1][4][ 32 ];
assign rho_out[2][0][ 52 ] = rho_in[2][0][ 49 ];
assign rho_out[2][1][ 52 ] = rho_in[2][1][ 42 ];
assign rho_out[2][2][ 52 ] = rho_in[2][2][ 9 ];
assign rho_out[2][3][ 52 ] = rho_in[2][3][ 27 ];
assign rho_out[2][4][ 52 ] = rho_in[2][4][ 13 ];
assign rho_out[3][0][ 52 ] = rho_in[3][0][ 11 ];
assign rho_out[3][1][ 52 ] = rho_in[3][1][ 7 ];
assign rho_out[3][2][ 52 ] = rho_in[3][2][ 37 ];
assign rho_out[3][3][ 52 ] = rho_in[3][3][ 31 ];
assign rho_out[3][4][ 52 ] = rho_in[3][4][ 44 ];
assign rho_out[4][0][ 52 ] = rho_in[4][0][ 34 ];
assign rho_out[4][1][ 52 ] = rho_in[4][1][ 50 ];
assign rho_out[4][2][ 52 ] = rho_in[4][2][ 55 ];
assign rho_out[4][3][ 52 ] = rho_in[4][3][ 60 ];
assign rho_out[4][4][ 52 ] = rho_in[4][4][ 38 ];
assign rho_out[0][0][ 53 ] = rho_in[0][0][ 53 ];
assign rho_out[0][1][ 53 ] = rho_in[0][1][ 52 ];
assign rho_out[0][2][ 53 ] = rho_in[0][2][ 55 ];
assign rho_out[0][3][ 53 ] = rho_in[0][3][ 25 ];
assign rho_out[0][4][ 53 ] = rho_in[0][4][ 26 ];
assign rho_out[1][0][ 53 ] = rho_in[1][0][ 17 ];
assign rho_out[1][1][ 53 ] = rho_in[1][1][ 9 ];
assign rho_out[1][2][ 53 ] = rho_in[1][2][ 47 ];
assign rho_out[1][3][ 53 ] = rho_in[1][3][ 62 ];
assign rho_out[1][4][ 53 ] = rho_in[1][4][ 33 ];
assign rho_out[2][0][ 53 ] = rho_in[2][0][ 50 ];
assign rho_out[2][1][ 53 ] = rho_in[2][1][ 43 ];
assign rho_out[2][2][ 53 ] = rho_in[2][2][ 10 ];
assign rho_out[2][3][ 53 ] = rho_in[2][3][ 28 ];
assign rho_out[2][4][ 53 ] = rho_in[2][4][ 14 ];
assign rho_out[3][0][ 53 ] = rho_in[3][0][ 12 ];
assign rho_out[3][1][ 53 ] = rho_in[3][1][ 8 ];
assign rho_out[3][2][ 53 ] = rho_in[3][2][ 38 ];
assign rho_out[3][3][ 53 ] = rho_in[3][3][ 32 ];
assign rho_out[3][4][ 53 ] = rho_in[3][4][ 45 ];
assign rho_out[4][0][ 53 ] = rho_in[4][0][ 35 ];
assign rho_out[4][1][ 53 ] = rho_in[4][1][ 51 ];
assign rho_out[4][2][ 53 ] = rho_in[4][2][ 56 ];
assign rho_out[4][3][ 53 ] = rho_in[4][3][ 61 ];
assign rho_out[4][4][ 53 ] = rho_in[4][4][ 39 ];
assign rho_out[0][0][ 54 ] = rho_in[0][0][ 54 ];
assign rho_out[0][1][ 54 ] = rho_in[0][1][ 53 ];
assign rho_out[0][2][ 54 ] = rho_in[0][2][ 56 ];
assign rho_out[0][3][ 54 ] = rho_in[0][3][ 26 ];
assign rho_out[0][4][ 54 ] = rho_in[0][4][ 27 ];
assign rho_out[1][0][ 54 ] = rho_in[1][0][ 18 ];
assign rho_out[1][1][ 54 ] = rho_in[1][1][ 10 ];
assign rho_out[1][2][ 54 ] = rho_in[1][2][ 48 ];
assign rho_out[1][3][ 54 ] = rho_in[1][3][ 63 ];
assign rho_out[1][4][ 54 ] = rho_in[1][4][ 34 ];
assign rho_out[2][0][ 54 ] = rho_in[2][0][ 51 ];
assign rho_out[2][1][ 54 ] = rho_in[2][1][ 44 ];
assign rho_out[2][2][ 54 ] = rho_in[2][2][ 11 ];
assign rho_out[2][3][ 54 ] = rho_in[2][3][ 29 ];
assign rho_out[2][4][ 54 ] = rho_in[2][4][ 15 ];
assign rho_out[3][0][ 54 ] = rho_in[3][0][ 13 ];
assign rho_out[3][1][ 54 ] = rho_in[3][1][ 9 ];
assign rho_out[3][2][ 54 ] = rho_in[3][2][ 39 ];
assign rho_out[3][3][ 54 ] = rho_in[3][3][ 33 ];
assign rho_out[3][4][ 54 ] = rho_in[3][4][ 46 ];
assign rho_out[4][0][ 54 ] = rho_in[4][0][ 36 ];
assign rho_out[4][1][ 54 ] = rho_in[4][1][ 52 ];
assign rho_out[4][2][ 54 ] = rho_in[4][2][ 57 ];
assign rho_out[4][3][ 54 ] = rho_in[4][3][ 62 ];
assign rho_out[4][4][ 54 ] = rho_in[4][4][ 40 ];
assign rho_out[0][0][ 55 ] = rho_in[0][0][ 55 ];
assign rho_out[0][1][ 55 ] = rho_in[0][1][ 54 ];
assign rho_out[0][2][ 55 ] = rho_in[0][2][ 57 ];
assign rho_out[0][3][ 55 ] = rho_in[0][3][ 27 ];
assign rho_out[0][4][ 55 ] = rho_in[0][4][ 28 ];
assign rho_out[1][0][ 55 ] = rho_in[1][0][ 19 ];
assign rho_out[1][1][ 55 ] = rho_in[1][1][ 11 ];
assign rho_out[1][2][ 55 ] = rho_in[1][2][ 49 ];
assign rho_out[1][3][ 55 ] = rho_in[1][3][ 0 ];
assign rho_out[1][4][ 55 ] = rho_in[1][4][ 35 ];
assign rho_out[2][0][ 55 ] = rho_in[2][0][ 52 ];
assign rho_out[2][1][ 55 ] = rho_in[2][1][ 45 ];
assign rho_out[2][2][ 55 ] = rho_in[2][2][ 12 ];
assign rho_out[2][3][ 55 ] = rho_in[2][3][ 30 ];
assign rho_out[2][4][ 55 ] = rho_in[2][4][ 16 ];
assign rho_out[3][0][ 55 ] = rho_in[3][0][ 14 ];
assign rho_out[3][1][ 55 ] = rho_in[3][1][ 10 ];
assign rho_out[3][2][ 55 ] = rho_in[3][2][ 40 ];
assign rho_out[3][3][ 55 ] = rho_in[3][3][ 34 ];
assign rho_out[3][4][ 55 ] = rho_in[3][4][ 47 ];
assign rho_out[4][0][ 55 ] = rho_in[4][0][ 37 ];
assign rho_out[4][1][ 55 ] = rho_in[4][1][ 53 ];
assign rho_out[4][2][ 55 ] = rho_in[4][2][ 58 ];
assign rho_out[4][3][ 55 ] = rho_in[4][3][ 63 ];
assign rho_out[4][4][ 55 ] = rho_in[4][4][ 41 ];
assign rho_out[0][0][ 56 ] = rho_in[0][0][ 56 ];
assign rho_out[0][1][ 56 ] = rho_in[0][1][ 55 ];
assign rho_out[0][2][ 56 ] = rho_in[0][2][ 58 ];
assign rho_out[0][3][ 56 ] = rho_in[0][3][ 28 ];
assign rho_out[0][4][ 56 ] = rho_in[0][4][ 29 ];
assign rho_out[1][0][ 56 ] = rho_in[1][0][ 20 ];
assign rho_out[1][1][ 56 ] = rho_in[1][1][ 12 ];
assign rho_out[1][2][ 56 ] = rho_in[1][2][ 50 ];
assign rho_out[1][3][ 56 ] = rho_in[1][3][ 1 ];
assign rho_out[1][4][ 56 ] = rho_in[1][4][ 36 ];
assign rho_out[2][0][ 56 ] = rho_in[2][0][ 53 ];
assign rho_out[2][1][ 56 ] = rho_in[2][1][ 46 ];
assign rho_out[2][2][ 56 ] = rho_in[2][2][ 13 ];
assign rho_out[2][3][ 56 ] = rho_in[2][3][ 31 ];
assign rho_out[2][4][ 56 ] = rho_in[2][4][ 17 ];
assign rho_out[3][0][ 56 ] = rho_in[3][0][ 15 ];
assign rho_out[3][1][ 56 ] = rho_in[3][1][ 11 ];
assign rho_out[3][2][ 56 ] = rho_in[3][2][ 41 ];
assign rho_out[3][3][ 56 ] = rho_in[3][3][ 35 ];
assign rho_out[3][4][ 56 ] = rho_in[3][4][ 48 ];
assign rho_out[4][0][ 56 ] = rho_in[4][0][ 38 ];
assign rho_out[4][1][ 56 ] = rho_in[4][1][ 54 ];
assign rho_out[4][2][ 56 ] = rho_in[4][2][ 59 ];
assign rho_out[4][3][ 56 ] = rho_in[4][3][ 0 ];
assign rho_out[4][4][ 56 ] = rho_in[4][4][ 42 ];
assign rho_out[0][0][ 57 ] = rho_in[0][0][ 57 ];
assign rho_out[0][1][ 57 ] = rho_in[0][1][ 56 ];
assign rho_out[0][2][ 57 ] = rho_in[0][2][ 59 ];
assign rho_out[0][3][ 57 ] = rho_in[0][3][ 29 ];
assign rho_out[0][4][ 57 ] = rho_in[0][4][ 30 ];
assign rho_out[1][0][ 57 ] = rho_in[1][0][ 21 ];
assign rho_out[1][1][ 57 ] = rho_in[1][1][ 13 ];
assign rho_out[1][2][ 57 ] = rho_in[1][2][ 51 ];
assign rho_out[1][3][ 57 ] = rho_in[1][3][ 2 ];
assign rho_out[1][4][ 57 ] = rho_in[1][4][ 37 ];
assign rho_out[2][0][ 57 ] = rho_in[2][0][ 54 ];
assign rho_out[2][1][ 57 ] = rho_in[2][1][ 47 ];
assign rho_out[2][2][ 57 ] = rho_in[2][2][ 14 ];
assign rho_out[2][3][ 57 ] = rho_in[2][3][ 32 ];
assign rho_out[2][4][ 57 ] = rho_in[2][4][ 18 ];
assign rho_out[3][0][ 57 ] = rho_in[3][0][ 16 ];
assign rho_out[3][1][ 57 ] = rho_in[3][1][ 12 ];
assign rho_out[3][2][ 57 ] = rho_in[3][2][ 42 ];
assign rho_out[3][3][ 57 ] = rho_in[3][3][ 36 ];
assign rho_out[3][4][ 57 ] = rho_in[3][4][ 49 ];
assign rho_out[4][0][ 57 ] = rho_in[4][0][ 39 ];
assign rho_out[4][1][ 57 ] = rho_in[4][1][ 55 ];
assign rho_out[4][2][ 57 ] = rho_in[4][2][ 60 ];
assign rho_out[4][3][ 57 ] = rho_in[4][3][ 1 ];
assign rho_out[4][4][ 57 ] = rho_in[4][4][ 43 ];
assign rho_out[0][0][ 58 ] = rho_in[0][0][ 58 ];
assign rho_out[0][1][ 58 ] = rho_in[0][1][ 57 ];
assign rho_out[0][2][ 58 ] = rho_in[0][2][ 60 ];
assign rho_out[0][3][ 58 ] = rho_in[0][3][ 30 ];
assign rho_out[0][4][ 58 ] = rho_in[0][4][ 31 ];
assign rho_out[1][0][ 58 ] = rho_in[1][0][ 22 ];
assign rho_out[1][1][ 58 ] = rho_in[1][1][ 14 ];
assign rho_out[1][2][ 58 ] = rho_in[1][2][ 52 ];
assign rho_out[1][3][ 58 ] = rho_in[1][3][ 3 ];
assign rho_out[1][4][ 58 ] = rho_in[1][4][ 38 ];
assign rho_out[2][0][ 58 ] = rho_in[2][0][ 55 ];
assign rho_out[2][1][ 58 ] = rho_in[2][1][ 48 ];
assign rho_out[2][2][ 58 ] = rho_in[2][2][ 15 ];
assign rho_out[2][3][ 58 ] = rho_in[2][3][ 33 ];
assign rho_out[2][4][ 58 ] = rho_in[2][4][ 19 ];
assign rho_out[3][0][ 58 ] = rho_in[3][0][ 17 ];
assign rho_out[3][1][ 58 ] = rho_in[3][1][ 13 ];
assign rho_out[3][2][ 58 ] = rho_in[3][2][ 43 ];
assign rho_out[3][3][ 58 ] = rho_in[3][3][ 37 ];
assign rho_out[3][4][ 58 ] = rho_in[3][4][ 50 ];
assign rho_out[4][0][ 58 ] = rho_in[4][0][ 40 ];
assign rho_out[4][1][ 58 ] = rho_in[4][1][ 56 ];
assign rho_out[4][2][ 58 ] = rho_in[4][2][ 61 ];
assign rho_out[4][3][ 58 ] = rho_in[4][3][ 2 ];
assign rho_out[4][4][ 58 ] = rho_in[4][4][ 44 ];
assign rho_out[0][0][ 59 ] = rho_in[0][0][ 59 ];
assign rho_out[0][1][ 59 ] = rho_in[0][1][ 58 ];
assign rho_out[0][2][ 59 ] = rho_in[0][2][ 61 ];
assign rho_out[0][3][ 59 ] = rho_in[0][3][ 31 ];
assign rho_out[0][4][ 59 ] = rho_in[0][4][ 32 ];
assign rho_out[1][0][ 59 ] = rho_in[1][0][ 23 ];
assign rho_out[1][1][ 59 ] = rho_in[1][1][ 15 ];
assign rho_out[1][2][ 59 ] = rho_in[1][2][ 53 ];
assign rho_out[1][3][ 59 ] = rho_in[1][3][ 4 ];
assign rho_out[1][4][ 59 ] = rho_in[1][4][ 39 ];
assign rho_out[2][0][ 59 ] = rho_in[2][0][ 56 ];
assign rho_out[2][1][ 59 ] = rho_in[2][1][ 49 ];
assign rho_out[2][2][ 59 ] = rho_in[2][2][ 16 ];
assign rho_out[2][3][ 59 ] = rho_in[2][3][ 34 ];
assign rho_out[2][4][ 59 ] = rho_in[2][4][ 20 ];
assign rho_out[3][0][ 59 ] = rho_in[3][0][ 18 ];
assign rho_out[3][1][ 59 ] = rho_in[3][1][ 14 ];
assign rho_out[3][2][ 59 ] = rho_in[3][2][ 44 ];
assign rho_out[3][3][ 59 ] = rho_in[3][3][ 38 ];
assign rho_out[3][4][ 59 ] = rho_in[3][4][ 51 ];
assign rho_out[4][0][ 59 ] = rho_in[4][0][ 41 ];
assign rho_out[4][1][ 59 ] = rho_in[4][1][ 57 ];
assign rho_out[4][2][ 59 ] = rho_in[4][2][ 62 ];
assign rho_out[4][3][ 59 ] = rho_in[4][3][ 3 ];
assign rho_out[4][4][ 59 ] = rho_in[4][4][ 45 ];
assign rho_out[0][0][ 60 ] = rho_in[0][0][ 60 ];
assign rho_out[0][1][ 60 ] = rho_in[0][1][ 59 ];
assign rho_out[0][2][ 60 ] = rho_in[0][2][ 62 ];
assign rho_out[0][3][ 60 ] = rho_in[0][3][ 32 ];
assign rho_out[0][4][ 60 ] = rho_in[0][4][ 33 ];
assign rho_out[1][0][ 60 ] = rho_in[1][0][ 24 ];
assign rho_out[1][1][ 60 ] = rho_in[1][1][ 16 ];
assign rho_out[1][2][ 60 ] = rho_in[1][2][ 54 ];
assign rho_out[1][3][ 60 ] = rho_in[1][3][ 5 ];
assign rho_out[1][4][ 60 ] = rho_in[1][4][ 40 ];
assign rho_out[2][0][ 60 ] = rho_in[2][0][ 57 ];
assign rho_out[2][1][ 60 ] = rho_in[2][1][ 50 ];
assign rho_out[2][2][ 60 ] = rho_in[2][2][ 17 ];
assign rho_out[2][3][ 60 ] = rho_in[2][3][ 35 ];
assign rho_out[2][4][ 60 ] = rho_in[2][4][ 21 ];
assign rho_out[3][0][ 60 ] = rho_in[3][0][ 19 ];
assign rho_out[3][1][ 60 ] = rho_in[3][1][ 15 ];
assign rho_out[3][2][ 60 ] = rho_in[3][2][ 45 ];
assign rho_out[3][3][ 60 ] = rho_in[3][3][ 39 ];
assign rho_out[3][4][ 60 ] = rho_in[3][4][ 52 ];
assign rho_out[4][0][ 60 ] = rho_in[4][0][ 42 ];
assign rho_out[4][1][ 60 ] = rho_in[4][1][ 58 ];
assign rho_out[4][2][ 60 ] = rho_in[4][2][ 63 ];
assign rho_out[4][3][ 60 ] = rho_in[4][3][ 4 ];
assign rho_out[4][4][ 60 ] = rho_in[4][4][ 46 ];
assign rho_out[0][0][ 61 ] = rho_in[0][0][ 61 ];
assign rho_out[0][1][ 61 ] = rho_in[0][1][ 60 ];
assign rho_out[0][2][ 61 ] = rho_in[0][2][ 63 ];
assign rho_out[0][3][ 61 ] = rho_in[0][3][ 33 ];
assign rho_out[0][4][ 61 ] = rho_in[0][4][ 34 ];
assign rho_out[1][0][ 61 ] = rho_in[1][0][ 25 ];
assign rho_out[1][1][ 61 ] = rho_in[1][1][ 17 ];
assign rho_out[1][2][ 61 ] = rho_in[1][2][ 55 ];
assign rho_out[1][3][ 61 ] = rho_in[1][3][ 6 ];
assign rho_out[1][4][ 61 ] = rho_in[1][4][ 41 ];
assign rho_out[2][0][ 61 ] = rho_in[2][0][ 58 ];
assign rho_out[2][1][ 61 ] = rho_in[2][1][ 51 ];
assign rho_out[2][2][ 61 ] = rho_in[2][2][ 18 ];
assign rho_out[2][3][ 61 ] = rho_in[2][3][ 36 ];
assign rho_out[2][4][ 61 ] = rho_in[2][4][ 22 ];
assign rho_out[3][0][ 61 ] = rho_in[3][0][ 20 ];
assign rho_out[3][1][ 61 ] = rho_in[3][1][ 16 ];
assign rho_out[3][2][ 61 ] = rho_in[3][2][ 46 ];
assign rho_out[3][3][ 61 ] = rho_in[3][3][ 40 ];
assign rho_out[3][4][ 61 ] = rho_in[3][4][ 53 ];
assign rho_out[4][0][ 61 ] = rho_in[4][0][ 43 ];
assign rho_out[4][1][ 61 ] = rho_in[4][1][ 59 ];
assign rho_out[4][2][ 61 ] = rho_in[4][2][ 0 ];
assign rho_out[4][3][ 61 ] = rho_in[4][3][ 5 ];
assign rho_out[4][4][ 61 ] = rho_in[4][4][ 47 ];
assign rho_out[0][0][ 62 ] = rho_in[0][0][ 62 ];
assign rho_out[0][1][ 62 ] = rho_in[0][1][ 61 ];
assign rho_out[0][2][ 62 ] = rho_in[0][2][ 0 ];
assign rho_out[0][3][ 62 ] = rho_in[0][3][ 34 ];
assign rho_out[0][4][ 62 ] = rho_in[0][4][ 35 ];
assign rho_out[1][0][ 62 ] = rho_in[1][0][ 26 ];
assign rho_out[1][1][ 62 ] = rho_in[1][1][ 18 ];
assign rho_out[1][2][ 62 ] = rho_in[1][2][ 56 ];
assign rho_out[1][3][ 62 ] = rho_in[1][3][ 7 ];
assign rho_out[1][4][ 62 ] = rho_in[1][4][ 42 ];
assign rho_out[2][0][ 62 ] = rho_in[2][0][ 59 ];
assign rho_out[2][1][ 62 ] = rho_in[2][1][ 52 ];
assign rho_out[2][2][ 62 ] = rho_in[2][2][ 19 ];
assign rho_out[2][3][ 62 ] = rho_in[2][3][ 37 ];
assign rho_out[2][4][ 62 ] = rho_in[2][4][ 23 ];
assign rho_out[3][0][ 62 ] = rho_in[3][0][ 21 ];
assign rho_out[3][1][ 62 ] = rho_in[3][1][ 17 ];
assign rho_out[3][2][ 62 ] = rho_in[3][2][ 47 ];
assign rho_out[3][3][ 62 ] = rho_in[3][3][ 41 ];
assign rho_out[3][4][ 62 ] = rho_in[3][4][ 54 ];
assign rho_out[4][0][ 62 ] = rho_in[4][0][ 44 ];
assign rho_out[4][1][ 62 ] = rho_in[4][1][ 60 ];
assign rho_out[4][2][ 62 ] = rho_in[4][2][ 1 ];
assign rho_out[4][3][ 62 ] = rho_in[4][3][ 6 ];
assign rho_out[4][4][ 62 ] = rho_in[4][4][ 48 ];
assign rho_out[0][0][ 63 ] = rho_in[0][0][ 63 ];
assign rho_out[0][1][ 63 ] = rho_in[0][1][ 62 ];
assign rho_out[0][2][ 63 ] = rho_in[0][2][ 1 ];
assign rho_out[0][3][ 63 ] = rho_in[0][3][ 35 ];
assign rho_out[0][4][ 63 ] = rho_in[0][4][ 36 ];
assign rho_out[1][0][ 63 ] = rho_in[1][0][ 27 ];
assign rho_out[1][1][ 63 ] = rho_in[1][1][ 19 ];
assign rho_out[1][2][ 63 ] = rho_in[1][2][ 57 ];
assign rho_out[1][3][ 63 ] = rho_in[1][3][ 8 ];
assign rho_out[1][4][ 63 ] = rho_in[1][4][ 43 ];
assign rho_out[2][0][ 63 ] = rho_in[2][0][ 60 ];
assign rho_out[2][1][ 63 ] = rho_in[2][1][ 53 ];
assign rho_out[2][2][ 63 ] = rho_in[2][2][ 20 ];
assign rho_out[2][3][ 63 ] = rho_in[2][3][ 38 ];
assign rho_out[2][4][ 63 ] = rho_in[2][4][ 24 ];
assign rho_out[3][0][ 63 ] = rho_in[3][0][ 22 ];
assign rho_out[3][1][ 63 ] = rho_in[3][1][ 18 ];
assign rho_out[3][2][ 63 ] = rho_in[3][2][ 48 ];
assign rho_out[3][3][ 63 ] = rho_in[3][3][ 42 ];
assign rho_out[3][4][ 63 ] = rho_in[3][4][ 55 ];
assign rho_out[4][0][ 63 ] = rho_in[4][0][ 45 ];
assign rho_out[4][1][ 63 ] = rho_in[4][1][ 61 ];
assign rho_out[4][2][ 63 ] = rho_in[4][2][ 2 ];
assign rho_out[4][3][ 63 ] = rho_in[4][3][ 7 ];
assign rho_out[4][4][ 63 ] = rho_in[4][4][ 49 ];


genvar hh;
generate
    for (hh = 0; hh <= N-1; hh = hh + 1) begin 
        assign iota_out[0][0][hh] = iota_in[0][0][hh] ^ Round_constant_signal[hh];
    end
endgenerate


function integer ABS;
    input integer numberIn;
    begin
        ABS = (numberIn < 0) ? -numberIn : numberIn;
    end
endfunction

endmodule
